module tg68k_alu_2_1_2_2
  (input  clk,
   input  reset,
   input  clkena_lw,
   input  [1:0] cpu,
   input  execopc,
   input  decodeopc,
   input  exe_condition,
   input  exec_tas,
   input  long_start,
   input  non_aligned,
   input  check_aligned,
   input  movem_presub,
   input  set_stop,
   input  z_error,
   input  [1:0] rot_bits,
   input  [88:0] exec,
   input  [31:0] op1out,
   input  [31:0] op2out,
   input  [31:0] reg_qa,
   input  [31:0] reg_qb,
   input  [15:0] opcode,
   input  [15:0] exe_opcode,
   input  [1:0] exe_datatype,
   input  [15:0] sndopc,
   input  [15:0] last_data_read,
   input  [15:0] data_read,
   input  [7:0] flagssr,
   input  [6:0] micro_state,
   input  [7:0] bf_ext_in,
   input  [5:0] bf_shift,
   input  [5:0] bf_width,
   input  [31:0] bf_ffo_offset,
   input  [4:0] bf_loffset,
   output [7:0] bf_ext_out,
   output set_v_flag,
   output [7:0] flags,
   output [2:0] c_out,
   output [31:0] addsub_q,
   output [31:0] aluout);
  wire [31:0] op1in;
  wire [31:0] addsub_a;
  wire [31:0] addsub_b;
  wire [33:0] notaddsub_b;
  wire [33:0] add_result;
  wire [2:0] addsub_ofl;
  wire opaddsub;
  wire [3:0] c_in;
  wire [2:0] flag_z;
  wire [3:0] set_flags;
  wire [7:0] ccrin;
  wire [3:0] last_flags1;
  wire [9:0] bcd_pur;
  wire [8:0] bcd_kor;
  wire halve_carry;
  wire vflag_a;
  wire bcd_a_carry;
  wire [8:0] bcd_a;
  wire [127:0] result_mulu;
  wire [63:0] result_div;
  wire [31:0] result_div_pre;
  wire set_mv_flag;
  wire v_flag;
  wire rot_rot;
  wire rot_x;
  wire rot_c;
  wire [31:0] rot_out;
  wire asl_vflag;
  wire [4:0] bit_number;
  wire [31:0] bits_out;
  wire one_bit_in;
  wire bchg;
  wire bset;
  wire [63:0] mulu_reg;
  wire [31:0] faktora;
  wire [31:0] faktorb;
  wire [63:0] div_reg;
  wire [63:0] div_quot;
  wire div_neg;
  wire div_bit;
  wire [32:0] div_sub;
  wire [32:0] div_over;
  wire nozero;
  wire div_qsign;
  wire [63:0] dividend;
  wire divs;
  wire signedop;
  wire op1_sign;
  wire [15:0] op2outext;
  wire [31:0] datareg;
  wire [31:0] bf_datareg;
  wire [39:0] result;
  wire [39:0] result_tmp;
  wire [31:0] unshifted_bitmask;
  wire [39:0] inmux0;
  wire [39:0] inmux1;
  wire [39:0] inmux2;
  wire [31:0] inmux3;
  wire [39:0] shifted_bitmask;
  wire [37:0] bitmaskmux0;
  wire [35:0] bitmaskmux1;
  wire [31:0] bitmaskmux2;
  wire [31:0] bitmaskmux3;
  wire [31:0] bf_set2;
  wire [39:0] shift;
  wire [5:0] bf_firstbit;
  wire [3:0] mux;
  wire [4:0] bitnr;
  wire [31:0] mask;
  wire mask_not_zero;
  wire bf_bset;
  wire bf_nflag;
  wire bf_bchg;
  wire bf_ins;
  wire bf_exts;
  wire bf_fffo;
  wire bf_d32;
  wire bf_s32;
  wire [33:0] hot_msb;
  wire [32:0] vector;
  wire [65:0] result_bs;
  wire [5:0] bit_nr;
  wire [5:0] bit_msb;
  wire [5:0] bs_shift;
  wire [5:0] bs_shift_mod;
  wire [32:0] asl_over;
  wire [32:0] asl_over_xor;
  wire [32:0] asr_sign;
  wire msb;
  wire [5:0] ring;
  wire [31:0] alu;
  wire [31:0] bsout;
  wire bs_v;
  wire bs_c;
  wire bs_x;
  wire n9439;
  wire n9440;
  wire [23:0] n9441;
  wire [6:0] n9442;
  wire n9443;
  wire [31:0] n9444;
  wire [31:0] n9445;
  wire [31:0] n9446;
  wire [31:0] n9447;
  wire [31:0] n9448;
  wire [31:0] n9449;
  wire n9450;
  wire n9451;
  wire n9452;
  wire [7:0] n9453;
  wire n9454;
  wire n9456;
  wire n9457;
  wire [31:0] n9458;
  wire [31:0] n9459;
  wire [31:0] n9460;
  wire n9461;
  wire n9463;
  wire n9464;
  wire n9466;
  wire [15:0] n9467;
  wire [15:0] n9468;
  wire [31:0] n9469;
  wire n9470;
  wire [31:0] n9471;
  wire [31:0] n9472;
  wire [31:0] n9473;
  wire [31:0] n9474;
  wire n9475;
  wire [31:0] n9476;
  wire n9477;
  wire [31:0] n9478;
  wire n9479;
  wire [3:0] n9480;
  wire [3:0] n9481;
  wire [7:0] n9482;
  wire n9483;
  wire [31:0] n9484;
  wire n9485;
  wire n9486;
  wire n9487;
  wire n9488;
  wire [15:0] n9489;
  wire [15:0] n9490;
  wire [31:0] n9491;
  wire n9492;
  wire n9493;
  wire n9494;
  wire n9495;
  wire [7:0] n9497;
  wire n9498;
  wire [3:0] n9499;
  wire [3:0] n9500;
  wire [7:0] n9501;
  wire [7:0] n9502;
  wire [7:0] n9503;
  wire [15:0] n9504;
  wire [7:0] n9505;
  wire [7:0] n9506;
  wire [7:0] n9507;
  wire [7:0] n9508;
  wire [7:0] n9509;
  wire [15:0] n9510;
  wire [15:0] n9511;
  wire [15:0] n9512;
  wire [15:0] n9513;
  wire [15:0] n9514;
  wire [15:0] n9515;
  wire [31:0] n9516;
  wire [31:0] n9517;
  wire [31:0] n9518;
  wire [31:0] n9519;
  wire [31:0] n9520;
  wire [31:0] n9521;
  wire [31:0] n9522;
  wire [7:0] n9523;
  wire [7:0] n9524;
  wire [23:0] n9525;
  wire [23:0] n9526;
  wire [23:0] n9527;
  wire [31:0] n9528;
  wire [31:0] n9529;
  wire [31:0] n9530;
  wire [31:0] n9531;
  wire [31:0] n9532;
  wire [7:0] n9533;
  wire [7:0] n9534;
  wire [23:0] n9535;
  wire [23:0] n9536;
  wire [23:0] n9537;
  wire n9542;
  wire n9543;
  wire n9544;
  wire n9545;
  wire [1:0] n9546;
  wire n9547;
  wire [2:0] n9548;
  wire [28:0] n9549;
  wire [31:0] n9550;
  wire [1:0] n9551;
  wire [31:0] n9553;
  wire [31:0] n9554;
  wire [31:0] n9555;
  wire n9556;
  wire n9559;
  wire n9561;
  wire [3:0] n9562;
  wire [7:0] n9564;
  wire [11:0] n9566;
  wire [3:0] n9567;
  wire [15:0] n9568;
  wire n9569;
  wire n9570;
  wire n9571;
  wire n9572;
  wire n9573;
  wire n9574;
  wire n9575;
  wire n9576;
  wire n9578;
  wire n9579;
  wire n9580;
  wire n9581;
  wire n9582;
  wire n9583;
  wire n9585;
  wire n9586;
  wire n9587;
  wire n9588;
  wire n9589;
  wire n9590;
  wire n9591;
  wire n9592;
  wire [31:0] n9595;
  wire [31:0] n9597;
  wire [31:0] n9599;
  wire n9600;
  wire n9601;
  wire n9602;
  wire n9603;
  wire n9604;
  wire n9606;
  wire n9607;
  wire [31:0] n9608;
  wire n9609;
  wire n9610;
  wire [15:0] n9611;
  wire [15:0] n9612;
  wire [15:0] n9613;
  wire [15:0] n9614;
  wire [15:0] n9615;
  wire n9617;
  wire n9618;
  wire n9619;
  wire n9620;
  wire n9621;
  wire n9622;
  wire n9623;
  wire [31:0] n9625;
  wire [31:0] n9626;
  wire n9627;
  wire n9628;
  wire n9630;
  wire [31:0] n9633;
  wire [31:0] n9634;
  wire [31:0] n9635;
  wire [31:0] n9636;
  wire [31:0] n9637;
  wire [31:0] n9638;
  wire n9639;
  wire n9640;
  wire [32:0] n9642;
  wire n9643;
  wire [33:0] n9644;
  wire [32:0] n9646;
  wire n9647;
  wire [33:0] n9648;
  wire [33:0] n9649;
  wire [33:0] n9650;
  wire [32:0] n9652;
  wire n9653;
  wire [33:0] n9654;
  wire [33:0] n9655;
  wire n9656;
  wire n9657;
  wire n9658;
  wire n9659;
  wire n9660;
  wire n9661;
  wire n9662;
  wire n9663;
  wire n9664;
  wire n9665;
  wire n9666;
  wire [31:0] n9667;
  wire n9668;
  wire n9669;
  wire n9670;
  wire n9671;
  wire n9672;
  wire n9673;
  wire n9674;
  wire n9675;
  wire n9676;
  wire n9677;
  wire n9678;
  wire n9679;
  wire n9680;
  wire n9681;
  wire n9682;
  wire n9683;
  wire n9684;
  wire n9685;
  wire n9686;
  wire n9687;
  wire n9688;
  wire [2:0] n9689;
  wire n9693;
  wire [8:0] n9694;
  wire [9:0] n9695;
  wire n9696;
  wire n9697;
  wire n9698;
  wire n9699;
  wire n9700;
  wire [3:0] n9703;
  localparam [8:0] n9704 = 9'b000000000;
  wire n9706;
  wire [3:0] n9708;
  wire [3:0] n9709;
  wire n9710;
  wire n9711;
  wire n9712;
  wire n9713;
  wire n9714;
  wire n9715;
  wire [8:0] n9716;
  wire [8:0] n9717;
  wire n9718;
  wire n9719;
  wire n9720;
  wire n9721;
  wire n9722;
  wire [3:0] n9724;
  wire n9725;
  wire n9726;
  wire n9727;
  wire n9728;
  wire n9729;
  wire n9730;
  wire n9731;
  wire n9732;
  wire n9733;
  wire n9734;
  wire n9735;
  wire n9736;
  wire n9737;
  wire [3:0] n9739;
  wire n9740;
  wire n9741;
  wire n9742;
  wire n9743;
  wire [8:0] n9744;
  wire [8:0] n9745;
  wire [7:0] n9746;
  wire [7:0] n9747;
  wire [7:0] n9748;
  wire n9749;
  wire [8:0] n9750;
  wire n9751;
  wire n9753;
  wire n9754;
  wire n9755;
  wire n9756;
  wire [1:0] n9761;
  wire n9763;
  wire n9765;
  wire [1:0] n9766;
  reg n9769;
  reg n9773;
  wire n9779;
  wire n9780;
  wire [1:0] n9781;
  wire n9783;
  wire [4:0] n9784;
  wire [2:0] n9785;
  wire [4:0] n9787;
  wire [4:0] n9788;
  wire [1:0] n9789;
  wire n9791;
  wire [4:0] n9792;
  wire [2:0] n9793;
  wire [4:0] n9795;
  wire [4:0] n9796;
  wire [4:0] n9797;
  wire n9803;
  wire n9804;
  wire n9805;
  wire [1:0] n9811;
  wire n9813;
  wire n9816;
  wire [2:0] n9818;
  wire n9820;
  wire n9822;
  wire n9824;
  wire n9826;
  wire n9828;
  wire [4:0] n9829;
  reg n9832;
  reg n9836;
  reg n9840;
  reg n9844;
  reg n9848;
  reg n9851;
  wire [1:0] n9852;
  wire n9854;
  wire n9857;
  wire [7:0] n9859;
  wire [31:0] n9876;
  wire [4:0] n9877;
  wire n9879;
  wire n9882;
  wire n9883;
  wire n9886;
  localparam [31:0] n9887 = 32'b00000000000000000000000000000000;
  wire [4:0] n9889;
  wire n9891;
  wire n9894;
  wire n9895;
  wire n9897;
  wire n9898;
  wire [4:0] n9900;
  wire n9902;
  wire n9905;
  wire n9906;
  wire n9908;
  wire n9909;
  wire [4:0] n9911;
  wire n9913;
  wire n9916;
  wire n9917;
  wire n9919;
  wire n9920;
  wire [4:0] n9922;
  wire n9924;
  wire n9927;
  wire n9928;
  wire n9930;
  wire n9931;
  wire [4:0] n9933;
  wire n9935;
  wire n9938;
  wire n9939;
  wire n9941;
  wire n9942;
  wire [4:0] n9944;
  wire n9946;
  wire n9949;
  wire n9950;
  wire n9952;
  wire n9953;
  wire [4:0] n9955;
  wire n9957;
  wire n9960;
  wire n9961;
  wire n9963;
  wire n9964;
  wire [4:0] n9966;
  wire n9968;
  wire n9971;
  wire n9972;
  wire n9974;
  wire n9975;
  wire [4:0] n9977;
  wire n9979;
  wire n9982;
  wire n9983;
  wire n9985;
  wire n9986;
  wire [4:0] n9988;
  wire n9990;
  wire n9993;
  wire n9994;
  wire n9996;
  wire n9997;
  wire [4:0] n9999;
  wire n10001;
  wire n10004;
  wire n10005;
  wire n10007;
  wire n10008;
  wire [4:0] n10010;
  wire n10012;
  wire n10015;
  wire n10016;
  wire n10018;
  wire n10019;
  wire [4:0] n10021;
  wire n10023;
  wire n10026;
  wire n10027;
  wire n10029;
  wire n10030;
  wire [4:0] n10032;
  wire n10034;
  wire n10037;
  wire n10038;
  wire n10040;
  wire n10041;
  wire [4:0] n10043;
  wire n10045;
  wire n10048;
  wire n10049;
  wire n10051;
  wire n10052;
  wire [4:0] n10054;
  wire n10056;
  wire n10059;
  wire n10060;
  wire n10062;
  wire n10063;
  wire [4:0] n10065;
  wire n10067;
  wire n10070;
  wire n10071;
  wire n10073;
  wire n10074;
  wire [4:0] n10076;
  wire n10078;
  wire n10081;
  wire n10082;
  wire n10084;
  wire n10085;
  wire [4:0] n10087;
  wire n10089;
  wire n10092;
  wire n10093;
  wire n10095;
  wire n10096;
  wire [4:0] n10098;
  wire n10100;
  wire n10103;
  wire n10104;
  wire n10106;
  wire n10107;
  wire [4:0] n10109;
  wire n10111;
  wire n10114;
  wire n10115;
  wire n10117;
  wire n10118;
  wire [4:0] n10120;
  wire n10122;
  wire n10125;
  wire n10126;
  wire n10128;
  wire n10129;
  wire [4:0] n10131;
  wire n10133;
  wire n10136;
  wire n10137;
  wire n10139;
  wire n10140;
  wire [4:0] n10142;
  wire n10144;
  wire n10147;
  wire n10148;
  wire n10150;
  wire n10151;
  wire [4:0] n10153;
  wire n10155;
  wire n10158;
  wire n10159;
  wire n10161;
  wire n10162;
  wire [4:0] n10164;
  wire n10166;
  wire n10169;
  wire n10170;
  wire n10172;
  wire n10173;
  wire [4:0] n10175;
  wire n10177;
  wire n10180;
  wire n10181;
  wire n10183;
  wire n10184;
  wire [4:0] n10186;
  wire n10188;
  wire n10191;
  wire n10192;
  wire n10194;
  wire n10195;
  wire [4:0] n10197;
  wire n10199;
  wire n10202;
  wire n10203;
  wire n10205;
  wire n10206;
  wire [4:0] n10208;
  wire n10210;
  wire n10213;
  wire n10214;
  wire n10215;
  wire n10216;
  wire n10217;
  wire n10218;
  wire [4:0] n10219;
  wire n10221;
  wire n10224;
  wire n10225;
  wire [4:0] n10227;
  wire n10230;
  wire [31:0] n10231;
  wire [31:0] n10232;
  wire n10233;
  wire [15:0] n10234;
  wire [15:0] n10235;
  wire [31:0] n10236;
  wire [31:0] n10237;
  wire n10238;
  wire [23:0] n10239;
  wire [7:0] n10240;
  wire [31:0] n10241;
  wire [31:0] n10242;
  wire n10243;
  wire [35:0] n10245;
  wire [3:0] n10246;
  wire [3:0] n10247;
  wire [3:0] n10248;
  wire [31:0] n10249;
  wire [35:0] n10251;
  wire [35:0] n10252;
  wire [35:0] n10253;
  wire n10254;
  wire [37:0] n10256;
  wire [1:0] n10257;
  wire [1:0] n10258;
  wire [1:0] n10259;
  wire [35:0] n10260;
  wire [37:0] n10262;
  wire [37:0] n10263;
  wire [37:0] n10264;
  wire n10265;
  wire [38:0] n10267;
  wire [39:0] n10269;
  wire n10270;
  wire n10271;
  wire n10272;
  wire [38:0] n10273;
  wire [39:0] n10275;
  wire [39:0] n10276;
  wire [39:0] n10277;
  wire [39:0] n10278;
  wire [7:0] n10279;
  wire [7:0] n10280;
  wire [7:0] n10281;
  wire [31:0] n10282;
  wire n10283;
  wire n10284;
  wire [38:0] n10285;
  wire [39:0] n10286;
  wire [39:0] n10287;
  wire n10288;
  wire [1:0] n10289;
  wire [37:0] n10290;
  wire [39:0] n10291;
  wire [39:0] n10292;
  wire n10293;
  wire [3:0] n10294;
  wire [35:0] n10295;
  wire [39:0] n10296;
  wire [39:0] n10297;
  wire n10298;
  wire [7:0] n10299;
  wire [23:0] n10300;
  wire [31:0] n10301;
  wire [31:0] n10302;
  wire [31:0] n10303;
  wire n10304;
  wire [15:0] n10305;
  wire [15:0] n10306;
  wire [31:0] n10307;
  wire [31:0] n10308;
  wire [7:0] n10309;
  wire [31:0] n10310;
  wire [7:0] n10311;
  wire [39:0] n10312;
  wire [39:0] n10314;
  wire [39:0] n10315;
  wire [39:0] n10316;
  wire [39:0] n10318;
  wire [39:0] n10319;
  wire [39:0] n10320;
  wire [39:0] n10321;
  wire n10322;
  wire n10323;
  wire n10324;
  wire n10325;
  wire n10327;
  wire n10328;
  wire n10329;
  wire n10330;
  wire n10332;
  wire n10333;
  wire n10334;
  wire n10335;
  wire n10337;
  wire n10338;
  wire n10339;
  wire n10340;
  wire n10342;
  wire n10343;
  wire n10344;
  wire n10345;
  wire n10347;
  wire n10348;
  wire n10349;
  wire n10350;
  wire n10352;
  wire n10353;
  wire n10354;
  wire n10355;
  wire n10357;
  wire n10358;
  wire n10359;
  wire n10360;
  wire n10362;
  wire n10363;
  wire n10364;
  wire n10365;
  wire n10367;
  wire n10368;
  wire n10369;
  wire n10370;
  wire n10372;
  wire n10373;
  wire n10374;
  wire n10375;
  wire n10377;
  wire n10378;
  wire n10379;
  wire n10380;
  wire n10382;
  wire n10383;
  wire n10384;
  wire n10385;
  wire n10387;
  wire n10388;
  wire n10389;
  wire n10390;
  wire n10392;
  wire n10393;
  wire n10394;
  wire n10395;
  wire n10397;
  wire n10398;
  wire n10399;
  wire n10400;
  wire n10402;
  wire n10403;
  wire n10404;
  wire n10405;
  wire n10407;
  wire n10408;
  wire n10409;
  wire n10410;
  wire n10412;
  wire n10413;
  wire n10414;
  wire n10415;
  wire n10417;
  wire n10418;
  wire n10419;
  wire n10420;
  wire n10422;
  wire n10423;
  wire n10424;
  wire n10425;
  wire n10427;
  wire n10428;
  wire n10429;
  wire n10430;
  wire n10432;
  wire n10433;
  wire n10434;
  wire n10435;
  wire n10437;
  wire n10438;
  wire n10439;
  wire n10440;
  wire n10442;
  wire n10443;
  wire n10444;
  wire n10445;
  wire n10447;
  wire n10448;
  wire n10449;
  wire n10450;
  wire n10452;
  wire n10453;
  wire n10454;
  wire n10455;
  wire n10457;
  wire n10458;
  wire n10459;
  wire n10460;
  wire n10462;
  wire n10463;
  wire n10464;
  wire n10465;
  wire n10467;
  wire n10468;
  wire n10469;
  wire n10470;
  wire n10472;
  wire n10473;
  wire n10474;
  wire n10475;
  wire n10477;
  wire n10478;
  wire n10479;
  wire n10480;
  wire n10482;
  wire n10483;
  wire n10484;
  wire n10485;
  wire n10487;
  wire n10488;
  wire n10489;
  wire n10490;
  wire n10492;
  wire n10493;
  wire n10494;
  wire n10495;
  wire n10497;
  wire n10498;
  wire n10499;
  wire n10500;
  wire n10502;
  wire n10503;
  wire n10504;
  wire n10505;
  wire n10507;
  wire n10508;
  wire n10509;
  wire n10510;
  wire n10512;
  wire n10513;
  wire n10514;
  wire n10515;
  wire n10516;
  wire n10517;
  wire n10518;
  wire n10519;
  wire [5:0] n10521;
  wire [5:0] n10522;
  wire [5:0] n10523;
  wire [3:0] n10524;
  wire n10526;
  wire [3:0] n10527;
  wire n10529;
  wire [3:0] n10530;
  wire n10532;
  wire [3:0] n10533;
  wire n10535;
  wire [3:0] n10537;
  wire n10539;
  wire [3:0] n10540;
  wire n10542;
  wire [3:0] n10544;
  wire n10546;
  wire [3:0] n10548;
  wire [3:0] n10549;
  wire [3:0] n10550;
  wire n10552;
  wire [3:0] n10553;
  wire [3:0] n10555;
  wire [1:0] n10556;
  wire n10557;
  wire n10558;
  wire n10559;
  wire n10561;
  wire [3:0] n10562;
  wire [3:0] n10563;
  wire [1:0] n10564;
  wire [1:0] n10566;
  wire [3:0] n10567;
  wire [3:0] n10570;
  wire [1:0] n10571;
  wire [2:0] n10572;
  wire [1:0] n10573;
  wire [1:0] n10574;
  wire n10575;
  wire n10577;
  wire [3:0] n10578;
  wire [3:0] n10580;
  wire [2:0] n10581;
  wire n10582;
  wire n10584;
  wire n10585;
  wire n10586;
  wire n10587;
  wire n10589;
  wire [3:0] n10590;
  wire [3:0] n10592;
  wire [2:0] n10593;
  wire n10594;
  wire n10595;
  wire [1:0] n10596;
  wire [1:0] n10598;
  wire [3:0] n10599;
  wire [3:0] n10600;
  wire [2:0] n10601;
  wire [2:0] n10603;
  localparam [4:0] n10604 = 5'b11111;
  wire [1:0] n10606;
  wire n10608;
  wire n10610;
  wire n10611;
  wire n10613;
  wire n10614;
  wire n10617;
  wire n10618;
  wire n10619;
  wire n10621;
  wire n10622;
  wire n10623;
  wire n10625;
  wire n10626;
  wire [1:0] n10627;
  wire n10628;
  wire n10629;
  wire n10630;
  wire n10631;
  wire n10632;
  wire n10635;
  wire [1:0] n10640;
  wire n10641;
  wire n10643;
  wire n10644;
  wire n10646;
  wire n10648;
  wire n10649;
  wire n10650;
  wire n10652;
  wire [2:0] n10653;
  reg n10654;
  wire n10672;
  wire n10673;
  wire n10675;
  wire n10676;
  wire n10678;
  wire n10679;
  wire n10682;
  wire n10683;
  wire n10703;
  wire n10704;
  wire n10707;
  wire n10708;
  wire [31:0] n10709;
  wire n10714;
  wire [1:0] n10715;
  wire n10717;
  wire n10719;
  wire n10721;
  wire n10722;
  wire n10724;
  wire [2:0] n10725;
  reg [5:0] n10730;
  wire [1:0] n10731;
  wire n10733;
  wire n10735;
  wire n10737;
  wire n10738;
  wire n10740;
  wire [2:0] n10741;
  reg [5:0] n10746;
  wire [5:0] n10747;
  wire [1:0] n10749;
  wire n10751;
  wire n10752;
  wire n10753;
  wire n10754;
  wire n10755;
  wire [5:0] n10756;
  wire [2:0] n10757;
  wire [2:0] n10758;
  wire n10760;
  wire [2:0] n10763;
  wire [5:0] n10764;
  wire [5:0] n10765;
  wire [5:0] n10767;
  localparam [33:0] n10770 = 34'b0000000000000000000000000000000000;
  wire n10774;
  wire [5:0] n10775;
  wire [5:0] n10777;
  wire [30:0] n10779;
  wire [31:0] n10781;
  wire [30:0] n10782;
  wire [31:0] n10784;
  wire [31:0] n10785;
  wire [32:0] n10786;
  wire [1:0] n10787;
  wire n10790;
  wire n10793;
  wire n10795;
  wire n10796;
  wire [1:0] n10797;
  wire n10798;
  reg n10799;
  wire n10800;
  reg n10801;
  wire [7:0] n10803;
  wire [15:0] n10804;
  wire [6:0] n10805;
  wire [31:0] n10806;
  wire [32:0] n10808;
  wire [32:0] n10809;
  wire n10811;
  wire n10812;
  wire n10813;
  wire n10814;
  wire n10815;
  wire n10817;
  wire n10819;
  wire n10820;
  wire n10821;
  wire [1:0] n10822;
  wire n10823;
  wire n10825;
  wire n10826;
  wire n10828;
  wire n10830;
  wire n10831;
  wire n10832;
  wire n10834;
  wire [2:0] n10835;
  reg n10836;
  wire n10837;
  wire n10839;
  wire n10840;
  wire [1:0] n10841;
  wire [7:0] n10842;
  wire [7:0] n10843;
  wire [7:0] n10844;
  wire n10845;
  wire n10847;
  wire [15:0] n10848;
  wire [15:0] n10849;
  wire [15:0] n10850;
  wire n10851;
  wire n10853;
  wire n10855;
  wire n10856;
  wire [31:0] n10857;
  wire [31:0] n10858;
  wire [31:0] n10859;
  wire n10860;
  wire n10862;
  wire [2:0] n10863;
  wire [7:0] n10864;
  wire [7:0] n10865;
  reg [7:0] n10867;
  wire [7:0] n10868;
  wire [7:0] n10869;
  reg [7:0] n10871;
  wire [15:0] n10872;
  reg [15:0] n10874;
  reg n10875;
  wire n10876;
  wire n10877;
  wire n10878;
  wire n10880;
  wire [1:0] n10881;
  wire [7:0] n10882;
  wire [7:0] n10883;
  wire [7:0] n10884;
  wire n10885;
  wire n10886;
  wire n10887;
  wire n10889;
  wire [15:0] n10890;
  wire [15:0] n10891;
  wire [15:0] n10892;
  wire n10893;
  wire n10894;
  wire n10895;
  wire n10897;
  wire n10899;
  wire n10900;
  wire [31:0] n10901;
  wire [31:0] n10902;
  wire [31:0] n10903;
  wire n10904;
  wire n10905;
  wire n10906;
  wire n10908;
  wire [2:0] n10909;
  wire [7:0] n10910;
  wire [7:0] n10911;
  reg [7:0] n10913;
  wire [7:0] n10914;
  wire [7:0] n10915;
  reg [7:0] n10917;
  wire [15:0] n10918;
  reg [15:0] n10920;
  reg n10921;
  wire n10922;
  wire n10923;
  wire [31:0] n10924;
  wire [31:0] n10925;
  wire [31:0] n10926;
  wire [31:0] n10927;
  wire [31:0] n10928;
  wire n10929;
  wire [31:0] n10930;
  wire [31:0] n10931;
  wire n10933;
  wire n10934;
  wire n10936;
  wire n10938;
  wire n10939;
  wire n10941;
  wire n10942;
  wire n10944;
  wire n10945;
  wire n10946;
  wire n10948;
  wire n10950;
  wire [5:0] n10952;
  wire n10954;
  wire [5:0] n10956;
  wire n10958;
  wire [5:0] n10960;
  wire n10962;
  wire [5:0] n10964;
  wire n10966;
  wire [5:0] n10968;
  wire n10970;
  wire [5:0] n10972;
  wire [5:0] n10973;
  wire [5:0] n10974;
  wire [5:0] n10975;
  wire [5:0] n10976;
  wire [5:0] n10977;
  wire [5:0] n10978;
  wire [5:0] n10980;
  wire n10982;
  wire n10984;
  wire [5:0] n10986;
  wire n10988;
  wire [5:0] n10990;
  wire n10992;
  wire [5:0] n10994;
  wire [5:0] n10995;
  wire [5:0] n10996;
  wire [5:0] n10997;
  wire n10999;
  wire n11001;
  wire [5:0] n11003;
  wire [5:0] n11004;
  wire n11006;
  wire [2:0] n11007;
  wire [5:0] n11009;
  wire n11011;
  wire [3:0] n11012;
  wire [5:0] n11014;
  wire n11016;
  wire [4:0] n11017;
  wire [5:0] n11019;
  wire n11021;
  wire [5:0] n11022;
  reg [5:0] n11024;
  wire n11025;
  wire n11026;
  wire [5:0] n11027;
  wire [5:0] n11028;
  wire n11029;
  wire n11030;
  wire n11031;
  wire n11032;
  wire [5:0] n11034;
  wire [5:0] n11035;
  wire n11036;
  wire n11037;
  wire n11038;
  wire [5:0] n11040;
  wire [5:0] n11041;
  wire [5:0] n11042;
  wire n11043;
  wire n11044;
  wire n11045;
  wire [5:0] n11047;
  wire [5:0] n11049;
  wire n11051;
  wire [5:0] n11052;
  wire n11053;
  wire [5:0] n11054;
  wire n11055;
  wire [31:0] n11056;
  wire [31:0] n11057;
  wire [31:0] n11058;
  localparam [32:0] n11059 = 33'b000000000000000000000000000000000;
  wire n11060;
  wire n11062;
  wire n11063;
  wire n11064;
  wire n11065;
  wire n11066;
  wire [31:0] n11067;
  wire [31:0] n11068;
  wire n11069;
  wire n11071;
  wire [31:0] n11072;
  wire n11073;
  wire [32:0] n11075;
  wire [1:0] n11076;
  wire n11077;
  localparam [23:0] n11078 = 24'b000000000000000000000000;
  localparam [23:0] n11079 = 24'b000000000000000000000000;
  wire n11081;
  wire n11082;
  wire n11083;
  wire n11084;
  wire [22:0] n11085;
  wire n11087;
  wire n11088;
  localparam [15:0] n11089 = 16'b0000000000000000;
  wire n11092;
  wire n11093;
  wire n11094;
  wire n11095;
  wire [14:0] n11096;
  wire n11098;
  wire n11100;
  wire n11101;
  wire n11102;
  wire n11104;
  wire n11105;
  wire n11106;
  wire n11107;
  wire n11109;
  wire [2:0] n11110;
  wire n11111;
  reg n11112;
  wire [6:0] n11113;
  wire [6:0] n11114;
  reg [6:0] n11115;
  wire n11116;
  wire n11117;
  reg n11118;
  wire [14:0] n11119;
  wire [14:0] n11120;
  reg [14:0] n11121;
  wire n11122;
  reg n11123;
  wire [7:0] n11125;
  reg n11129;
  wire [7:0] n11130;
  wire [7:0] n11131;
  reg [7:0] n11132;
  wire [15:0] n11133;
  wire [15:0] n11134;
  reg [15:0] n11135;
  wire [7:0] n11137;
  wire [65:0] n11139;
  wire [30:0] n11140;
  wire [31:0] n11141;
  wire [65:0] n11142;
  wire n11146;
  wire [7:0] n11147;
  wire [7:0] n11148;
  wire n11149;
  wire [7:0] n11150;
  wire [7:0] n11151;
  wire n11152;
  wire [7:0] n11153;
  wire [7:0] n11154;
  wire [7:0] n11155;
  wire [7:0] n11156;
  wire [7:0] n11157;
  wire [7:0] n11158;
  wire n11159;
  wire n11160;
  wire n11161;
  wire n11162;
  wire [7:0] n11163;
  wire n11165;
  wire [7:0] n11167;
  wire n11169;
  wire [15:0] n11171;
  wire n11173;
  wire n11176;
  wire [1:0] n11177;
  wire [1:0] n11179;
  wire [2:0] n11180;
  wire [2:0] n11182;
  wire [2:0] n11184;
  wire n11187;
  wire n11188;
  wire n11189;
  wire [1:0] n11190;
  wire n11191;
  wire [2:0] n11192;
  wire n11193;
  wire [3:0] n11194;
  wire n11195;
  wire n11196;
  wire n11197;
  wire [1:0] n11198;
  wire [1:0] n11199;
  wire [1:0] n11200;
  wire [1:0] n11201;
  wire n11203;
  wire n11204;
  wire n11205;
  wire n11206;
  wire n11207;
  wire [1:0] n11208;
  wire n11209;
  wire [2:0] n11210;
  wire n11211;
  wire [3:0] n11212;
  wire n11213;
  wire n11214;
  wire [1:0] n11215;
  wire n11216;
  wire [2:0] n11217;
  wire n11218;
  wire [3:0] n11219;
  wire [3:0] n11220;
  wire [3:0] n11221;
  wire [3:0] n11222;
  wire n11224;
  wire n11225;
  wire [7:0] n11226;
  wire [7:0] n11227;
  wire n11228;
  wire [7:0] n11229;
  wire [7:0] n11230;
  wire n11231;
  wire n11232;
  wire n11233;
  wire n11234;
  wire n11235;
  wire n11236;
  wire n11238;
  wire n11239;
  wire n11241;
  wire n11242;
  wire n11243;
  wire n11244;
  wire n11245;
  wire [1:0] n11247;
  wire [3:0] n11249;
  wire [3:0] n11251;
  wire [3:0] n11252;
  wire [3:0] n11253;
  wire n11254;
  wire n11255;
  wire [3:0] n11256;
  wire n11257;
  wire n11258;
  wire n11259;
  wire n11261;
  wire n11262;
  wire n11263;
  wire n11264;
  wire n11265;
  wire n11266;
  wire n11267;
  wire n11268;
  wire n11269;
  wire n11270;
  wire n11271;
  wire n11272;
  wire n11273;
  wire n11274;
  wire n11276;
  wire n11278;
  wire n11280;
  wire n11281;
  wire n11282;
  wire [1:0] n11283;
  wire [3:0] n11285;
  wire n11286;
  wire n11287;
  wire [1:0] n11288;
  wire [3:0] n11290;
  wire [3:0] n11291;
  wire [3:0] n11292;
  wire n11293;
  wire n11295;
  wire n11296;
  wire n11297;
  wire n11298;
  wire n11299;
  wire n11302;
  wire n11304;
  wire n11305;
  wire n11306;
  wire n11308;
  wire n11309;
  wire n11310;
  wire n11311;
  wire n11312;
  wire n11313;
  wire n11314;
  wire n11315;
  wire n11316;
  wire n11317;
  wire n11318;
  wire n11319;
  wire n11320;
  wire n11321;
  wire n11323;
  wire n11324;
  wire n11327;
  wire n11328;
  wire n11329;
  wire n11330;
  wire n11331;
  wire [1:0] n11332;
  wire n11334;
  wire n11335;
  wire n11336;
  wire n11337;
  wire n11338;
  wire n11341;
  wire n11342;
  wire [1:0] n11343;
  wire n11344;
  wire n11345;
  wire n11346;
  wire n11347;
  wire n11348;
  wire n11349;
  wire n11350;
  wire n11351;
  wire n11352;
  wire n11353;
  wire n11354;
  wire n11355;
  wire n11356;
  wire n11357;
  wire n11358;
  wire n11359;
  wire n11360;
  wire n11361;
  wire n11362;
  wire n11363;
  wire n11364;
  wire n11365;
  wire n11367;
  wire n11368;
  wire n11369;
  wire n11370;
  wire n11371;
  wire n11372;
  wire n11374;
  wire n11375;
  wire n11376;
  wire n11377;
  wire [15:0] n11378;
  wire n11380;
  wire n11382;
  wire [15:0] n11383;
  wire n11385;
  wire n11386;
  wire n11387;
  wire n11390;
  wire [3:0] n11393;
  wire [3:0] n11394;
  wire [3:0] n11395;
  wire [3:0] n11396;
  wire [3:0] n11397;
  wire [1:0] n11398;
  wire [1:0] n11399;
  wire [1:0] n11400;
  wire n11401;
  wire n11402;
  wire n11403;
  wire n11404;
  wire n11405;
  wire [3:0] n11406;
  wire [3:0] n11407;
  wire [3:0] n11408;
  wire [3:0] n11409;
  wire [3:0] n11410;
  wire [3:0] n11411;
  wire [3:0] n11412;
  wire [3:0] n11413;
  wire [3:0] n11414;
  wire [3:0] n11415;
  wire [3:0] n11416;
  wire [3:0] n11417;
  wire [3:0] n11418;
  wire [4:0] n11419;
  wire [4:0] n11420;
  wire [4:0] n11421;
  wire [3:0] n11422;
  wire [3:0] n11423;
  wire [3:0] n11424;
  wire n11425;
  wire n11426;
  wire n11427;
  wire [3:0] n11428;
  wire [4:0] n11429;
  wire [4:0] n11430;
  wire [4:0] n11431;
  wire [2:0] n11432;
  wire [2:0] n11433;
  wire [2:0] n11434;
  wire [3:0] n11436;
  wire [7:0] n11437;
  wire [7:0] n11438;
  wire [3:0] n11439;
  wire n11440;
  wire [7:0] n11442;
  wire [3:0] n11443;
  wire n11444;
  wire [4:0] n11446;
  wire [7:0] n11447;
  wire n11454;
  wire n11455;
  wire n11456;
  wire [31:0] n11459;
  wire n11460;
  wire n11461;
  wire [31:0] n11464;
  wire [15:0] n11465;
  wire [15:0] n11466;
  wire n11467;
  wire n11468;
  wire [15:0] n11471;
  wire n11472;
  wire n11473;
  wire [15:0] n11476;
  wire [31:0] n11477;
  wire [31:0] n11478;
  wire [31:0] n11479;
  wire [31:0] n11480;
  wire [15:0] n11481;
  wire [47:0] n11482;
  wire [15:0] n11483;
  wire [63:0] n11484;
  wire [15:0] n11485;
  wire [47:0] n11486;
  wire [15:0] n11487;
  wire [63:0] n11488;
  wire [127:0] n11489;
  wire [127:0] n11490;
  wire [127:0] n11491;
  wire [31:0] n11492;
  wire n11494;
  wire n11495;
  wire n11496;
  wire n11497;
  wire n11498;
  wire n11499;
  wire [31:0] n11500;
  wire n11502;
  wire n11503;
  wire n11504;
  wire n11505;
  wire n11506;
  wire n11509;
  wire [31:0] n11514;
  wire n11522;
  wire n11523;
  wire n11524;
  wire n11525;
  wire n11526;
  wire n11527;
  wire n11528;
  wire n11529;
  wire n11531;
  wire n11532;
  wire n11533;
  wire n11534;
  wire n11535;
  wire n11536;
  wire n11537;
  wire n11538;
  wire n11539;
  wire n11540;
  wire n11541;
  wire n11542;
  wire n11543;
  wire n11544;
  wire n11545;
  wire n11546;
  wire n11547;
  wire n11548;
  wire n11549;
  wire n11550;
  wire n11551;
  wire n11552;
  wire n11553;
  wire n11554;
  wire n11555;
  wire n11556;
  wire n11557;
  wire n11558;
  wire n11559;
  wire n11560;
  wire n11561;
  wire n11562;
  wire n11563;
  wire n11564;
  wire n11565;
  wire n11566;
  wire n11567;
  wire n11568;
  wire n11569;
  wire n11570;
  wire n11571;
  wire n11572;
  wire n11573;
  wire n11574;
  wire n11575;
  wire n11576;
  wire n11577;
  wire n11578;
  wire n11579;
  wire n11580;
  wire n11581;
  wire n11582;
  wire n11583;
  wire n11584;
  wire n11585;
  wire n11586;
  wire n11587;
  wire n11588;
  wire n11589;
  wire n11590;
  wire n11591;
  wire n11592;
  wire n11593;
  wire n11594;
  wire [3:0] n11595;
  wire [3:0] n11596;
  wire [3:0] n11597;
  wire [3:0] n11598;
  wire [3:0] n11599;
  wire [3:0] n11600;
  wire [3:0] n11601;
  wire [3:0] n11602;
  wire [15:0] n11603;
  wire [15:0] n11604;
  wire [31:0] n11605;
  wire n11606;
  wire n11608;
  wire n11609;
  wire n11610;
  wire n11611;
  wire n11612;
  wire [31:0] n11613;
  wire n11614;
  wire n11615;
  wire [63:0] n11616;
  wire [15:0] n11617;
  wire [15:0] n11618;
  wire [31:0] n11619;
  wire [31:0] n11620;
  wire [15:0] n11621;
  wire [15:0] n11622;
  wire [15:0] n11623;
  wire n11625;
  wire n11626;
  wire n11627;
  wire [15:0] n11628;
  wire [15:0] n11630;
  wire n11631;
  wire n11632;
  wire [32:0] n11633;
  wire [32:0] n11635;
  wire [32:0] n11636;
  wire [32:0] n11637;
  wire [16:0] n11639;
  wire [15:0] n11640;
  wire [32:0] n11641;
  wire [32:0] n11642;
  wire [32:0] n11643;
  wire n11644;
  wire [31:0] n11645;
  wire [31:0] n11646;
  wire [31:0] n11647;
  wire [30:0] n11648;
  wire n11649;
  wire [31:0] n11650;
  wire [31:0] n11651;
  wire [31:0] n11653;
  wire [31:0] n11654;
  wire [31:0] n11655;
  wire n11656;
  wire n11657;
  wire n11658;
  wire n11659;
  wire n11660;
  wire n11661;
  wire n11662;
  wire n11663;
  wire n11664;
  wire n11665;
  wire n11666;
  wire n11667;
  wire n11669;
  wire n11672;
  wire n11678;
  wire n11681;
  wire n11682;
  wire n11683;
  wire [63:0] n11685;
  wire [63:0] n11686;
  wire n11689;
  wire n11690;
  wire n11691;
  wire [63:0] n11692;
  wire n11694;
  wire n11697;
  wire n11698;
  wire n11699;
  wire n11700;
  wire [31:0] n11701;
  wire [32:0] n11703;
  wire [16:0] n11705;
  wire [15:0] n11706;
  wire [32:0] n11707;
  wire [32:0] n11708;
  wire n11711;
  wire n11712;
  wire [31:0] n11713;
  wire [31:0] n11715;
  wire [31:0] n11716;
  wire [31:0] n11717;
  wire [63:0] n11718;
  wire n11720;
  wire n11721;
  wire n11723;
  wire n11724;
  wire n11727;
  wire [31:0] n11737;
  wire [2:0] n11738;
  wire [3:0] n11739;
  reg [3:0] n11740;
  wire [8:0] n11741;
  wire [63:0] n11742;
  reg [63:0] n11743;
  wire n11744;
  reg n11745;
  reg n11746;
  wire n11748;
  reg n11749;
  wire n11750;
  reg n11751;
  wire [31:0] n11755;
  wire [31:0] n11756;
  reg [31:0] n11757;
  wire [63:0] n11759;
  wire [63:0] n11761;
  reg [63:0] n11762;
  wire [63:0] n11763;
  wire n11765;
  reg n11766;
  wire [32:0] n11767;
  reg [32:0] n11768;
  wire n11769;
  reg n11770;
  wire [63:0] n11771;
  wire n11772;
  reg n11773;
  wire n11774;
  reg n11775;
  wire [31:0] n11778;
  wire [39:0] n11780;
  wire [31:0] n11781;
  wire [39:0] n11783;
  wire [4:0] n11784;
  wire n11785;
  reg n11786;
  wire n11787;
  reg n11788;
  wire n11789;
  reg n11790;
  wire n11791;
  reg n11792;
  wire n11793;
  reg n11794;
  wire n11795;
  reg n11796;
  wire n11797;
  reg n11798;
  wire [32:0] n11800;
  wire [32:0] n11801;
  wire [32:0] n11802;
  wire [31:0] n11803;
  wire [7:0] n11804;
  reg [7:0] n11805;
  reg [7:0] n11806;
  wire n11807;
  wire n11808;
  wire n11809;
  wire n11810;
  wire n11811;
  wire n11812;
  wire n11813;
  wire n11814;
  wire n11815;
  wire n11816;
  wire n11817;
  wire n11818;
  wire n11819;
  wire n11820;
  wire n11821;
  wire n11822;
  wire n11823;
  wire n11824;
  wire n11825;
  wire n11826;
  wire n11827;
  wire n11828;
  wire n11829;
  wire n11830;
  wire n11831;
  wire n11832;
  wire n11833;
  wire n11834;
  wire n11835;
  wire n11836;
  wire n11837;
  wire n11838;
  wire n11839;
  wire n11840;
  wire n11841;
  wire n11842;
  wire n11843;
  wire n11844;
  wire n11845;
  wire n11846;
  wire n11847;
  wire n11848;
  wire n11849;
  wire n11850;
  wire n11851;
  wire n11852;
  wire n11853;
  wire n11854;
  wire n11855;
  wire n11856;
  wire n11857;
  wire n11858;
  wire n11859;
  wire n11860;
  wire n11861;
  wire n11862;
  wire n11863;
  wire n11864;
  wire n11865;
  wire n11866;
  wire n11867;
  wire n11868;
  wire n11869;
  wire n11870;
  wire n11871;
  wire n11872;
  wire n11873;
  wire n11874;
  wire n11875;
  wire n11876;
  wire n11877;
  wire n11878;
  wire n11879;
  wire n11880;
  wire n11881;
  wire n11882;
  wire n11883;
  wire n11884;
  wire n11885;
  wire n11886;
  wire n11887;
  wire n11888;
  wire n11889;
  wire n11890;
  wire n11891;
  wire n11892;
  wire n11893;
  wire n11894;
  wire n11895;
  wire n11896;
  wire n11897;
  wire n11898;
  wire n11899;
  wire n11900;
  wire n11901;
  wire n11902;
  wire n11903;
  wire n11904;
  wire n11905;
  wire n11906;
  wire n11907;
  wire n11908;
  wire n11909;
  wire n11910;
  wire n11911;
  wire n11912;
  wire n11913;
  wire n11914;
  wire n11915;
  wire n11916;
  wire n11917;
  wire n11918;
  wire n11919;
  wire n11920;
  wire n11921;
  wire n11922;
  wire n11923;
  wire n11924;
  wire n11925;
  wire n11926;
  wire n11927;
  wire n11928;
  wire n11929;
  wire n11930;
  wire n11931;
  wire n11932;
  wire n11933;
  wire n11934;
  wire n11935;
  wire n11936;
  wire n11937;
  wire n11938;
  wire n11939;
  wire n11940;
  wire n11941;
  wire [31:0] n11942;
  wire n11943;
  wire n11944;
  wire n11945;
  wire n11946;
  wire n11947;
  wire n11948;
  wire n11949;
  wire n11950;
  wire n11951;
  wire n11952;
  wire n11953;
  wire n11954;
  wire n11955;
  wire n11956;
  wire n11957;
  wire n11958;
  wire n11959;
  wire n11960;
  wire n11961;
  wire n11962;
  wire n11963;
  wire n11964;
  wire n11965;
  wire n11966;
  wire n11967;
  wire n11968;
  wire n11969;
  wire n11970;
  wire n11971;
  wire n11972;
  wire n11973;
  wire n11974;
  wire n11975;
  wire n11976;
  wire n11977;
  wire n11978;
  wire n11979;
  wire n11980;
  wire n11981;
  wire n11982;
  wire n11983;
  wire n11984;
  wire n11985;
  wire n11986;
  wire n11987;
  wire n11988;
  wire n11989;
  wire n11990;
  wire n11991;
  wire n11992;
  wire n11993;
  wire n11994;
  wire n11995;
  wire n11996;
  wire n11997;
  wire n11998;
  wire n11999;
  wire n12000;
  wire n12001;
  wire n12002;
  wire n12003;
  wire n12004;
  wire n12005;
  wire n12006;
  wire n12007;
  wire n12008;
  wire n12009;
  wire n12010;
  wire n12011;
  wire n12012;
  wire n12013;
  wire n12014;
  wire n12015;
  wire n12016;
  wire n12017;
  wire n12018;
  wire n12019;
  wire n12020;
  wire n12021;
  wire n12022;
  wire n12023;
  wire n12024;
  wire n12025;
  wire n12026;
  wire n12027;
  wire n12028;
  wire n12029;
  wire n12030;
  wire n12031;
  wire n12032;
  wire n12033;
  wire n12034;
  wire n12035;
  wire n12036;
  wire n12037;
  wire n12038;
  wire n12039;
  wire n12040;
  wire n12041;
  wire n12042;
  wire n12043;
  wire n12044;
  wire n12045;
  wire n12046;
  wire n12047;
  wire n12048;
  wire n12049;
  wire n12050;
  wire n12051;
  wire n12052;
  wire n12053;
  wire n12054;
  wire n12055;
  wire n12056;
  wire n12057;
  wire n12058;
  wire n12059;
  wire n12060;
  wire n12061;
  wire n12062;
  wire n12063;
  wire n12064;
  wire n12065;
  wire n12066;
  wire n12067;
  wire n12068;
  wire n12069;
  wire n12070;
  wire n12071;
  wire n12072;
  wire n12073;
  wire n12074;
  wire n12075;
  wire n12076;
  wire n12077;
  wire n12078;
  wire n12079;
  wire n12080;
  wire n12081;
  wire n12082;
  wire n12083;
  wire n12084;
  wire n12085;
  wire n12086;
  wire n12087;
  wire n12088;
  wire n12089;
  wire n12090;
  wire n12091;
  wire [33:0] n12092;
  assign bf_ext_out = n11805; //(module output)
  assign set_v_flag = n11672; //(module output)
  assign flags = n11806; //(module output)
  assign c_out = n9689; //(module output)
  assign addsub_q = n9667; //(module output)
  assign aluout = n9449; //(module output)
  /* TG68K_ALU.vhd:86:16  */
  assign op1in = n11737; // (signal)
  /* TG68K_ALU.vhd:87:16  */
  assign addsub_a = n9555; // (signal)
  /* TG68K_ALU.vhd:88:16  */
  assign addsub_b = n9638; // (signal)
  /* TG68K_ALU.vhd:89:16  */
  assign notaddsub_b = n9650; // (signal)
  /* TG68K_ALU.vhd:90:16  */
  assign add_result = n9655; // (signal)
  /* TG68K_ALU.vhd:91:16  */
  assign addsub_ofl = n11738; // (signal)
  /* TG68K_ALU.vhd:92:16  */
  assign opaddsub = n9617; // (signal)
  /* TG68K_ALU.vhd:93:16  */
  assign c_in = n11739; // (signal)
  /* TG68K_ALU.vhd:94:16  */
  assign flag_z = n11184; // (signal)
  /* TG68K_ALU.vhd:95:16  */
  assign set_flags = n11222; // (signal)
  /* TG68K_ALU.vhd:96:16  */
  assign ccrin = n11158; // (signal)
  /* TG68K_ALU.vhd:97:16  */
  assign last_flags1 = n11740; // (signal)
  /* TG68K_ALU.vhd:100:16  */
  assign bcd_pur = n9695; // (signal)
  /* TG68K_ALU.vhd:101:16  */
  assign bcd_kor = n11741; // (signal)
  /* TG68K_ALU.vhd:102:16  */
  assign halve_carry = n9700; // (signal)
  /* TG68K_ALU.vhd:103:16  */
  assign vflag_a = n9753; // (signal)
  /* TG68K_ALU.vhd:104:16  */
  assign bcd_a_carry = n9756; // (signal)
  /* TG68K_ALU.vhd:105:16  */
  assign bcd_a = n9750; // (signal)
  /* TG68K_ALU.vhd:106:16  */
  assign result_mulu = n11491; // (signal)
  /* TG68K_ALU.vhd:107:16  */
  assign result_div = n11743; // (signal)
  /* TG68K_ALU.vhd:108:16  */
  assign result_div_pre = n11655; // (signal)
  /* TG68K_ALU.vhd:109:16  */
  assign set_mv_flag = n11509; // (signal)
  /* TG68K_ALU.vhd:110:16  */
  assign v_flag = n11745; // (signal)
  /* TG68K_ALU.vhd:112:16  */
  assign rot_rot = n10654; // (signal)
  /* TG68K_ALU.vhd:115:16  */
  assign rot_x = n10707; // (signal)
  /* TG68K_ALU.vhd:116:16  */
  assign rot_c = n10708; // (signal)
  /* TG68K_ALU.vhd:117:16  */
  assign rot_out = n10709; // (signal)
  /* TG68K_ALU.vhd:118:16  */
  assign asl_vflag = n11746; // (signal)
  /* TG68K_ALU.vhd:120:16  */
  assign bit_number = n9797; // (signal)
  /* TG68K_ALU.vhd:121:16  */
  assign bits_out = n11942; // (signal)
  /* TG68K_ALU.vhd:122:16  */
  assign one_bit_in = n11807; // (signal)
  /* TG68K_ALU.vhd:123:16  */
  assign bchg = n11749; // (signal)
  /* TG68K_ALU.vhd:124:16  */
  assign bset = n11751; // (signal)
  /* TG68K_ALU.vhd:129:16  */
  assign mulu_reg = n11759; // (signal)
  /* TG68K_ALU.vhd:131:16  */
  assign faktora = n11478; // (signal)
  /* TG68K_ALU.vhd:132:16  */
  assign faktorb = n11480; // (signal)
  /* TG68K_ALU.vhd:134:16  */
  assign div_reg = n11762; // (signal)
  /* TG68K_ALU.vhd:135:16  */
  assign div_quot = n11763; // (signal)
  /* TG68K_ALU.vhd:137:16  */
  assign div_neg = n11766; // (signal)
  /* TG68K_ALU.vhd:138:16  */
  assign div_bit = n11644; // (signal)
  /* TG68K_ALU.vhd:139:16  */
  assign div_sub = n11643; // (signal)
  /* TG68K_ALU.vhd:140:16  */
  assign div_over = n11768; // (signal)
  /* TG68K_ALU.vhd:141:16  */
  assign nozero = n11770; // (signal)
  /* TG68K_ALU.vhd:142:16  */
  assign div_qsign = n11615; // (signal)
  /* TG68K_ALU.vhd:143:16  */
  assign dividend = n11771; // (signal)
  /* TG68K_ALU.vhd:144:16  */
  assign divs = n11529; // (signal)
  /* TG68K_ALU.vhd:145:16  */
  assign signedop = n11773; // (signal)
  /* TG68K_ALU.vhd:146:16  */
  assign op1_sign = n11775; // (signal)
  /* TG68K_ALU.vhd:148:16  */
  assign op2outext = n11630; // (signal)
  /* TG68K_ALU.vhd:151:16  */
  assign datareg = n11778; // (signal)
  /* TG68K_ALU.vhd:153:16  */
  assign bf_datareg = n10232; // (signal)
  /* TG68K_ALU.vhd:154:16  */
  assign result = n11780; // (signal)
  /* TG68K_ALU.vhd:155:16  */
  assign result_tmp = n10321; // (signal)
  /* TG68K_ALU.vhd:156:16  */
  assign unshifted_bitmask = n11781; // (signal)
  /* TG68K_ALU.vhd:158:16  */
  assign inmux0 = n10287; // (signal)
  /* TG68K_ALU.vhd:159:16  */
  assign inmux1 = n10292; // (signal)
  /* TG68K_ALU.vhd:160:16  */
  assign inmux2 = n10297; // (signal)
  /* TG68K_ALU.vhd:161:16  */
  assign inmux3 = n10303; // (signal)
  /* TG68K_ALU.vhd:162:16  */
  assign shifted_bitmask = n10277; // (signal)
  /* TG68K_ALU.vhd:163:16  */
  assign bitmaskmux0 = n10264; // (signal)
  /* TG68K_ALU.vhd:164:16  */
  assign bitmaskmux1 = n10253; // (signal)
  /* TG68K_ALU.vhd:165:16  */
  assign bitmaskmux2 = n10242; // (signal)
  /* TG68K_ALU.vhd:166:16  */
  assign bitmaskmux3 = n10237; // (signal)
  /* TG68K_ALU.vhd:167:16  */
  assign bf_set2 = n10308; // (signal)
  /* TG68K_ALU.vhd:168:16  */
  assign shift = n11783; // (signal)
  /* TG68K_ALU.vhd:169:16  */
  assign bf_firstbit = n10523; // (signal)
  /* TG68K_ALU.vhd:170:16  */
  assign mux = n10600; // (signal)
  /* TG68K_ALU.vhd:171:16  */
  assign bitnr = n11784; // (signal)
  /* TG68K_ALU.vhd:172:16  */
  assign mask = datareg; // (signal)
  /* TG68K_ALU.vhd:173:16  */
  assign mask_not_zero = n10635; // (signal)
  /* TG68K_ALU.vhd:174:16  */
  assign bf_bset = n11786; // (signal)
  /* TG68K_ALU.vhd:175:16  */
  assign bf_nflag = n11943; // (signal)
  /* TG68K_ALU.vhd:176:16  */
  assign bf_bchg = n11788; // (signal)
  /* TG68K_ALU.vhd:177:16  */
  assign bf_ins = n11790; // (signal)
  /* TG68K_ALU.vhd:178:16  */
  assign bf_exts = n11792; // (signal)
  /* TG68K_ALU.vhd:179:16  */
  assign bf_fffo = n11794; // (signal)
  /* TG68K_ALU.vhd:180:16  */
  assign bf_d32 = n11796; // (signal)
  /* TG68K_ALU.vhd:181:16  */
  assign bf_s32 = n11798; // (signal)
  /* TG68K_ALU.vhd:187:16  */
  assign hot_msb = n12092; // (signal)
  /* TG68K_ALU.vhd:188:16  */
  assign vector = n11800; // (signal)
  /* TG68K_ALU.vhd:189:16  */
  assign result_bs = n11142; // (signal)
  /* TG68K_ALU.vhd:190:16  */
  assign bit_nr = n11054; // (signal)
  /* TG68K_ALU.vhd:191:16  */
  assign bit_msb = n10777; // (signal)
  /* TG68K_ALU.vhd:192:16  */
  assign bs_shift = n10767; // (signal)
  /* TG68K_ALU.vhd:193:16  */
  assign bs_shift_mod = n11024; // (signal)
  /* TG68K_ALU.vhd:194:16  */
  assign asl_over = n10809; // (signal)
  /* TG68K_ALU.vhd:195:16  */
  assign asl_over_xor = n11801; // (signal)
  /* TG68K_ALU.vhd:196:16  */
  assign asr_sign = n11802; // (signal)
  /* TG68K_ALU.vhd:197:16  */
  assign msb = n11129; // (signal)
  /* TG68K_ALU.vhd:198:16  */
  assign ring = n10747; // (signal)
  /* TG68K_ALU.vhd:199:16  */
  assign alu = n10931; // (signal)
  /* TG68K_ALU.vhd:200:16  */
  assign bsout = n11803; // (signal)
  /* TG68K_ALU.vhd:201:16  */
  assign bs_v = n10944; // (signal)
  /* TG68K_ALU.vhd:202:16  */
  assign bs_c = n11071; // (signal)
  /* TG68K_ALU.vhd:203:16  */
  assign bs_x = n10946; // (signal)
  /* TG68K_ALU.vhd:215:35  */
  assign n9439 = op1in[7]; // extract
  /* TG68K_ALU.vhd:215:39  */
  assign n9440 = n9439 | exec_tas;
  assign n9441 = op1in[31:8]; // extract
  assign n9442 = op1in[6:0]; // extract
  /* TG68K_ALU.vhd:216:24  */
  assign n9443 = exec[76]; // extract
  /* TG68K_ALU.vhd:217:41  */
  assign n9444 = result[31:0]; // extract
  /* TG68K_ALU.vhd:219:57  */
  assign n9445 = {26'b0, bf_firstbit};  //  uext
  /* TG68K_ALU.vhd:219:57  */
  assign n9446 = bf_ffo_offset - n9445;
  /* TG68K_ALU.vhd:218:25  */
  assign n9447 = bf_fffo ? n9446 : n9444;
  assign n9448 = {n9441, n9440, n9442};
  /* TG68K_ALU.vhd:216:17  */
  assign n9449 = n9443 ? n9447 : n9448;
  /* TG68K_ALU.vhd:224:24  */
  assign n9450 = exec[12]; // extract
  /* TG68K_ALU.vhd:224:45  */
  assign n9451 = exec[13]; // extract
  /* TG68K_ALU.vhd:224:38  */
  assign n9452 = n9450 | n9451;
  /* TG68K_ALU.vhd:225:51  */
  assign n9453 = bcd_a[7:0]; // extract
  /* TG68K_ALU.vhd:226:27  */
  assign n9454 = exec[20]; // extract
  /* TG68K_ALU.vhd:226:41  */
  assign n9456 = 1'b1 & n9454;
  /* TG68K_ALU.vhd:234:40  */
  assign n9457 = exec[67]; // extract
  /* TG68K_ALU.vhd:235:61  */
  assign n9458 = result_mulu[31:0]; // extract
  /* TG68K_ALU.vhd:238:58  */
  assign n9459 = mulu_reg[31:0]; // extract
  /* TG68K_ALU.vhd:234:33  */
  assign n9460 = n9457 ? n9458 : n9459;
  /* TG68K_ALU.vhd:241:27  */
  assign n9461 = exec[21]; // extract
  /* TG68K_ALU.vhd:241:41  */
  assign n9463 = 1'b1 & n9461;
  /* TG68K_ALU.vhd:242:38  */
  assign n9464 = exe_opcode[15]; // extract
  /* TG68K_ALU.vhd:242:47  */
  assign n9466 = n9464 | 1'b0;
  /* TG68K_ALU.vhd:244:52  */
  assign n9467 = result_div[47:32]; // extract
  /* TG68K_ALU.vhd:244:77  */
  assign n9468 = result_div[15:0]; // extract
  /* TG68K_ALU.vhd:244:66  */
  assign n9469 = {n9467, n9468};
  /* TG68K_ALU.vhd:246:40  */
  assign n9470 = exec[68]; // extract
  /* TG68K_ALU.vhd:247:60  */
  assign n9471 = result_div[63:32]; // extract
  /* TG68K_ALU.vhd:249:60  */
  assign n9472 = result_div[31:0]; // extract
  /* TG68K_ALU.vhd:246:33  */
  assign n9473 = n9470 ? n9471 : n9472;
  /* TG68K_ALU.vhd:242:25  */
  assign n9474 = n9466 ? n9469 : n9473;
  /* TG68K_ALU.vhd:252:27  */
  assign n9475 = exec[5]; // extract
  /* TG68K_ALU.vhd:253:41  */
  assign n9476 = op2out | op1out;
  /* TG68K_ALU.vhd:254:27  */
  assign n9477 = exec[6]; // extract
  /* TG68K_ALU.vhd:255:41  */
  assign n9478 = op2out & op1out;
  /* TG68K_ALU.vhd:256:27  */
  assign n9479 = exec[16]; // extract
  assign n9480 = {exe_condition, exe_condition, exe_condition, exe_condition};
  assign n9481 = {exe_condition, exe_condition, exe_condition, exe_condition};
  assign n9482 = {n9480, n9481};
  /* TG68K_ALU.vhd:258:27  */
  assign n9483 = exec[7]; // extract
  /* TG68K_ALU.vhd:259:41  */
  assign n9484 = op2out ^ op1out;
  /* TG68K_ALU.vhd:261:27  */
  assign n9485 = exec[85]; // extract
  /* TG68K_ALU.vhd:264:27  */
  assign n9486 = exec[9]; // extract
  /* TG68K_ALU.vhd:266:27  */
  assign n9487 = exec[81]; // extract
  /* TG68K_ALU.vhd:268:27  */
  assign n9488 = exec[15]; // extract
  /* TG68K_ALU.vhd:269:40  */
  assign n9489 = op1out[15:0]; // extract
  /* TG68K_ALU.vhd:269:61  */
  assign n9490 = op1out[31:16]; // extract
  /* TG68K_ALU.vhd:269:53  */
  assign n9491 = {n9489, n9490};
  /* TG68K_ALU.vhd:270:27  */
  assign n9492 = exec[14]; // extract
  /* TG68K_ALU.vhd:272:27  */
  assign n9493 = exec[75]; // extract
  /* TG68K_ALU.vhd:274:27  */
  assign n9494 = exec[2]; // extract
  /* TG68K_ALU.vhd:276:38  */
  assign n9495 = exe_opcode[9]; // extract
  /* TG68K_ALU.vhd:276:25  */
  assign n9497 = n9495 ? 8'b00000000 : flagssr;
  /* TG68K_ALU.vhd:281:27  */
  assign n9498 = exec[77]; // extract
  /* TG68K_ALU.vhd:282:54  */
  assign n9499 = n9667[11:8]; // extract
  /* TG68K_ALU.vhd:282:78  */
  assign n9500 = n9667[3:0]; // extract
  /* TG68K_ALU.vhd:282:68  */
  assign n9501 = {n9499, n9500};
  assign n9502 = n9667[7:0]; // extract
  /* TG68K_ALU.vhd:281:17  */
  assign n9503 = n9498 ? n9501 : n9502;
  assign n9504 = {n9497, n11806};
  assign n9505 = n9504[7:0]; // extract
  /* TG68K_ALU.vhd:274:17  */
  assign n9506 = n9494 ? n9505 : n9503;
  assign n9507 = n9504[15:8]; // extract
  assign n9508 = n9667[15:8]; // extract
  /* TG68K_ALU.vhd:274:17  */
  assign n9509 = n9494 ? n9507 : n9508;
  assign n9510 = {n9509, n9506};
  assign n9511 = bf_datareg[15:0]; // extract
  /* TG68K_ALU.vhd:272:17  */
  assign n9512 = n9493 ? n9511 : n9510;
  assign n9513 = bf_datareg[31:16]; // extract
  assign n9514 = n9667[31:16]; // extract
  /* TG68K_ALU.vhd:272:17  */
  assign n9515 = n9493 ? n9513 : n9514;
  assign n9516 = {n9515, n9512};
  /* TG68K_ALU.vhd:270:17  */
  assign n9517 = n9492 ? bits_out : n9516;
  /* TG68K_ALU.vhd:268:17  */
  assign n9518 = n9488 ? n9491 : n9517;
  /* TG68K_ALU.vhd:266:17  */
  assign n9519 = n9487 ? bsout : n9518;
  /* TG68K_ALU.vhd:264:17  */
  assign n9520 = n9486 ? rot_out : n9519;
  /* TG68K_ALU.vhd:261:17  */
  assign n9521 = n9485 ? op2out : n9520;
  /* TG68K_ALU.vhd:258:17  */
  assign n9522 = n9483 ? n9484 : n9521;
  assign n9523 = n9522[7:0]; // extract
  /* TG68K_ALU.vhd:256:17  */
  assign n9524 = n9479 ? n9482 : n9523;
  assign n9525 = n9522[31:8]; // extract
  assign n9526 = n9667[31:8]; // extract
  /* TG68K_ALU.vhd:256:17  */
  assign n9527 = n9479 ? n9526 : n9525;
  assign n9528 = {n9527, n9524};
  /* TG68K_ALU.vhd:254:17  */
  assign n9529 = n9477 ? n9478 : n9528;
  /* TG68K_ALU.vhd:252:17  */
  assign n9530 = n9475 ? n9476 : n9529;
  /* TG68K_ALU.vhd:241:17  */
  assign n9531 = n9463 ? n9474 : n9530;
  /* TG68K_ALU.vhd:226:17  */
  assign n9532 = n9456 ? n9460 : n9531;
  assign n9533 = n9532[7:0]; // extract
  /* TG68K_ALU.vhd:224:17  */
  assign n9534 = n9452 ? n9453 : n9533;
  assign n9535 = n9532[31:8]; // extract
  assign n9536 = n9667[31:8]; // extract
  /* TG68K_ALU.vhd:224:17  */
  assign n9537 = n9452 ? n9536 : n9535;
  /* TG68K_ALU.vhd:293:24  */
  assign n9542 = exec[29]; // extract
  /* TG68K_ALU.vhd:294:34  */
  assign n9543 = sndopc[11]; // extract
  /* TG68K_ALU.vhd:295:51  */
  assign n9544 = op1out[31]; // extract
  /* TG68K_ALU.vhd:295:62  */
  assign n9545 = op1out[31]; // extract
  /* TG68K_ALU.vhd:295:55  */
  assign n9546 = {n9544, n9545};
  /* TG68K_ALU.vhd:295:73  */
  assign n9547 = op1out[31]; // extract
  /* TG68K_ALU.vhd:295:66  */
  assign n9548 = {n9546, n9547};
  /* TG68K_ALU.vhd:295:84  */
  assign n9549 = op1out[31:3]; // extract
  /* TG68K_ALU.vhd:295:77  */
  assign n9550 = {n9548, n9549};
  /* TG68K_ALU.vhd:297:84  */
  assign n9551 = sndopc[10:9]; // extract
  /* TG68K_ALU.vhd:297:77  */
  assign n9553 = {30'b000000000000000000000000000000, n9551};
  /* TG68K_ALU.vhd:294:25  */
  assign n9554 = n9543 ? n9550 : n9553;
  /* TG68K_ALU.vhd:293:17  */
  assign n9555 = n9542 ? n9554 : op1out;
  /* TG68K_ALU.vhd:301:24  */
  assign n9556 = exec[48]; // extract
  /* TG68K_ALU.vhd:301:17  */
  assign n9559 = n9556 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:309:24  */
  assign n9561 = exec[78]; // extract
  /* TG68K_ALU.vhd:310:65  */
  assign n9562 = op2out[7:4]; // extract
  /* TG68K_ALU.vhd:310:57  */
  assign n9564 = {4'b0000, n9562};
  /* TG68K_ALU.vhd:310:78  */
  assign n9566 = {n9564, 4'b0000};
  /* TG68K_ALU.vhd:310:95  */
  assign n9567 = op2out[3:0]; // extract
  /* TG68K_ALU.vhd:310:87  */
  assign n9568 = {n9566, n9567};
  /* TG68K_ALU.vhd:311:30  */
  assign n9569 = ~execopc;
  /* TG68K_ALU.vhd:311:43  */
  assign n9570 = exec[53]; // extract
  /* TG68K_ALU.vhd:311:55  */
  assign n9571 = ~n9570;
  /* TG68K_ALU.vhd:311:35  */
  assign n9572 = n9571 & n9569;
  /* TG68K_ALU.vhd:311:68  */
  assign n9573 = exec[29]; // extract
  /* TG68K_ALU.vhd:311:82  */
  assign n9574 = ~n9573;
  /* TG68K_ALU.vhd:311:60  */
  assign n9575 = n9574 & n9572;
  /* TG68K_ALU.vhd:312:38  */
  assign n9576 = ~long_start;
  /* TG68K_ALU.vhd:312:59  */
  assign n9578 = exe_datatype == 2'b00;
  /* TG68K_ALU.vhd:312:43  */
  assign n9579 = n9578 & n9576;
  /* TG68K_ALU.vhd:312:73  */
  assign n9580 = exec[50]; // extract
  /* TG68K_ALU.vhd:312:81  */
  assign n9581 = ~n9580;
  /* TG68K_ALU.vhd:312:65  */
  assign n9582 = n9581 & n9579;
  /* TG68K_ALU.vhd:314:41  */
  assign n9583 = ~long_start;
  /* TG68K_ALU.vhd:314:62  */
  assign n9585 = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:314:46  */
  assign n9586 = n9585 & n9583;
  /* TG68K_ALU.vhd:314:77  */
  assign n9587 = exec[47]; // extract
  /* TG68K_ALU.vhd:314:93  */
  assign n9588 = exec[46]; // extract
  /* TG68K_ALU.vhd:314:86  */
  assign n9589 = n9587 | n9588;
  /* TG68K_ALU.vhd:314:103  */
  assign n9590 = n9589 | movem_presub;
  /* TG68K_ALU.vhd:314:68  */
  assign n9591 = n9590 & n9586;
  /* TG68K_ALU.vhd:315:40  */
  assign n9592 = exec[69]; // extract
  /* TG68K_ALU.vhd:315:33  */
  assign n9595 = n9592 ? 32'b00000000000000000000000000000110 : 32'b00000000000000000000000000000100;
  /* TG68K_ALU.vhd:314:25  */
  assign n9597 = n9591 ? n9595 : 32'b00000000000000000000000000000010;
  /* TG68K_ALU.vhd:312:25  */
  assign n9599 = n9582 ? 32'b00000000000000000000000000000001 : n9597;
  /* TG68K_ALU.vhd:324:33  */
  assign n9600 = exec[28]; // extract
  /* TG68K_ALU.vhd:324:59  */
  assign n9601 = n11806[4]; // extract
  /* TG68K_ALU.vhd:324:50  */
  assign n9602 = n9601 & n9600;
  /* TG68K_ALU.vhd:324:75  */
  assign n9603 = exec[31]; // extract
  /* TG68K_ALU.vhd:324:68  */
  assign n9604 = n9602 | n9603;
  /* TG68K_ALU.vhd:324:25  */
  assign n9606 = n9604 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:327:41  */
  assign n9607 = exec[56]; // extract
  /* TG68K_ALU.vhd:311:17  */
  assign n9608 = n9575 ? n9599 : op2out;
  /* TG68K_ALU.vhd:311:17  */
  assign n9609 = n9575 ? n9559 : n9607;
  /* TG68K_ALU.vhd:311:17  */
  assign n9610 = n9575 ? 1'b0 : n9606;
  /* TG68KdotC_Kernel.vhd:1283:1  */
  assign n9611 = n9608[15:0]; // extract
  /* TG68K_ALU.vhd:309:17  */
  assign n9612 = n9561 ? n9568 : n9611;
  /* TG68KdotC_Kernel.vhd:1254:17  */
  assign n9613 = n9608[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:1254:17  */
  assign n9614 = op2out[31:16]; // extract
  /* TG68K_ALU.vhd:309:17  */
  assign n9615 = n9561 ? n9614 : n9613;
  /* TG68K_ALU.vhd:309:17  */
  assign n9617 = n9561 ? n9559 : n9609;
  /* TG68K_ALU.vhd:309:17  */
  assign n9618 = n9561 ? 1'b0 : n9610;
  /* TG68K_ALU.vhd:331:24  */
  assign n9619 = exec[69]; // extract
  /* TG68K_ALU.vhd:331:43  */
  assign n9620 = n9619 | check_aligned;
  /* TG68K_ALU.vhd:332:36  */
  assign n9621 = ~movem_presub;
  /* TG68K_ALU.vhd:333:64  */
  assign n9622 = ~long_start;
  /* TG68K_ALU.vhd:333:48  */
  assign n9623 = n9622 & non_aligned;
  assign n9625 = {n9615, n9612};
  /* TG68K_ALU.vhd:333:25  */
  assign n9626 = n9623 ? 32'b00000000000000000000000000000000 : n9625;
  /* TG68K_ALU.vhd:337:64  */
  assign n9627 = ~long_start;
  /* TG68K_ALU.vhd:337:48  */
  assign n9628 = n9627 & non_aligned;
  /* TG68K_ALU.vhd:338:44  */
  assign n9630 = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:338:27  */
  assign n9633 = n9630 ? 32'b00000000000000000000000000001000 : 32'b00000000000000000000000000000100;
  /* TG68KdotC_Kernel.vhd:941:17  */
  assign n9634 = {n9615, n9612};
  /* TG68K_ALU.vhd:337:25  */
  assign n9635 = n9628 ? n9633 : n9634;
  /* TG68K_ALU.vhd:332:19  */
  assign n9636 = n9621 ? n9626 : n9635;
  /* TG68KdotC_Kernel.vhd:870:17  */
  assign n9637 = {n9615, n9612};
  /* TG68K_ALU.vhd:331:17  */
  assign n9638 = n9620 ? n9636 : n9637;
  /* TG68K_ALU.vhd:347:28  */
  assign n9639 = ~opaddsub;
  /* TG68K_ALU.vhd:347:33  */
  assign n9640 = n9639 | long_start;
  /* TG68K_ALU.vhd:348:43  */
  assign n9642 = {1'b0, addsub_b};
  /* TG68K_ALU.vhd:348:57  */
  assign n9643 = c_in[0]; // extract
  /* TG68K_ALU.vhd:348:52  */
  assign n9644 = {n9642, n9643};
  /* TG68K_ALU.vhd:350:48  */
  assign n9646 = {1'b0, addsub_b};
  /* TG68K_ALU.vhd:350:62  */
  assign n9647 = c_in[0]; // extract
  /* TG68K_ALU.vhd:350:57  */
  assign n9648 = {n9646, n9647};
  /* TG68K_ALU.vhd:350:40  */
  assign n9649 = ~n9648;
  /* TG68K_ALU.vhd:347:17  */
  assign n9650 = n9640 ? n9644 : n9649;
  /* TG68K_ALU.vhd:352:36  */
  assign n9652 = {1'b0, addsub_a};
  /* TG68K_ALU.vhd:352:57  */
  assign n9653 = notaddsub_b[0]; // extract
  /* TG68K_ALU.vhd:352:45  */
  assign n9654 = {n9652, n9653};
  /* TG68K_ALU.vhd:352:61  */
  assign n9655 = n9654 + notaddsub_b;
  /* TG68K_ALU.vhd:353:38  */
  assign n9656 = add_result[9]; // extract
  /* TG68K_ALU.vhd:353:54  */
  assign n9657 = addsub_a[8]; // extract
  /* TG68K_ALU.vhd:353:42  */
  assign n9658 = n9656 ^ n9657;
  /* TG68K_ALU.vhd:353:70  */
  assign n9659 = addsub_b[8]; // extract
  /* TG68K_ALU.vhd:353:58  */
  assign n9660 = n9658 ^ n9659;
  /* TG68K_ALU.vhd:354:38  */
  assign n9661 = add_result[17]; // extract
  /* TG68K_ALU.vhd:354:55  */
  assign n9662 = addsub_a[16]; // extract
  /* TG68K_ALU.vhd:354:43  */
  assign n9663 = n9661 ^ n9662;
  /* TG68K_ALU.vhd:354:72  */
  assign n9664 = addsub_b[16]; // extract
  /* TG68K_ALU.vhd:354:60  */
  assign n9665 = n9663 ^ n9664;
  /* TG68K_ALU.vhd:355:38  */
  assign n9666 = add_result[33]; // extract
  /* TG68K_ALU.vhd:356:39  */
  assign n9667 = add_result[32:1]; // extract
  /* TG68K_ALU.vhd:357:39  */
  assign n9668 = c_in[1]; // extract
  /* TG68K_ALU.vhd:357:57  */
  assign n9669 = add_result[8]; // extract
  /* TG68K_ALU.vhd:357:43  */
  assign n9670 = n9668 ^ n9669;
  /* TG68K_ALU.vhd:357:73  */
  assign n9671 = addsub_a[7]; // extract
  /* TG68K_ALU.vhd:357:61  */
  assign n9672 = n9670 ^ n9671;
  /* TG68K_ALU.vhd:357:89  */
  assign n9673 = addsub_b[7]; // extract
  /* TG68K_ALU.vhd:357:77  */
  assign n9674 = n9672 ^ n9673;
  /* TG68K_ALU.vhd:358:39  */
  assign n9675 = c_in[2]; // extract
  /* TG68K_ALU.vhd:358:57  */
  assign n9676 = add_result[16]; // extract
  /* TG68K_ALU.vhd:358:43  */
  assign n9677 = n9675 ^ n9676;
  /* TG68K_ALU.vhd:358:74  */
  assign n9678 = addsub_a[15]; // extract
  /* TG68K_ALU.vhd:358:62  */
  assign n9679 = n9677 ^ n9678;
  /* TG68K_ALU.vhd:358:91  */
  assign n9680 = addsub_b[15]; // extract
  /* TG68K_ALU.vhd:358:79  */
  assign n9681 = n9679 ^ n9680;
  /* TG68K_ALU.vhd:359:39  */
  assign n9682 = c_in[3]; // extract
  /* TG68K_ALU.vhd:359:57  */
  assign n9683 = add_result[32]; // extract
  /* TG68K_ALU.vhd:359:43  */
  assign n9684 = n9682 ^ n9683;
  /* TG68K_ALU.vhd:359:74  */
  assign n9685 = addsub_a[31]; // extract
  /* TG68K_ALU.vhd:359:62  */
  assign n9686 = n9684 ^ n9685;
  /* TG68K_ALU.vhd:359:91  */
  assign n9687 = addsub_b[31]; // extract
  /* TG68K_ALU.vhd:359:79  */
  assign n9688 = n9686 ^ n9687;
  /* TG68K_ALU.vhd:360:30  */
  assign n9689 = c_in[3:1]; // extract
  /* TG68K_ALU.vhd:370:32  */
  assign n9693 = c_in[1]; // extract
  /* TG68K_ALU.vhd:370:46  */
  assign n9694 = add_result[8:0]; // extract
  /* TG68K_ALU.vhd:370:35  */
  assign n9695 = {n9693, n9694};
  /* TG68K_ALU.vhd:372:38  */
  assign n9696 = op1out[4]; // extract
  /* TG68K_ALU.vhd:372:52  */
  assign n9697 = op2out[4]; // extract
  /* TG68K_ALU.vhd:372:42  */
  assign n9698 = n9696 ^ n9697;
  /* TG68K_ALU.vhd:372:67  */
  assign n9699 = bcd_pur[5]; // extract
  /* TG68K_ALU.vhd:372:56  */
  assign n9700 = n9698 ^ n9699;
  /* TG68K_ALU.vhd:373:17  */
  assign n9703 = halve_carry ? 4'b0110 : 4'b0000;
  /* TG68K_ALU.vhd:376:27  */
  assign n9706 = bcd_pur[9]; // extract
  assign n9708 = n9704[7:4]; // extract
  /* TG68K_ALU.vhd:376:17  */
  assign n9709 = n9706 ? 4'b0110 : n9708;
  assign n9710 = n9704[8]; // extract
  /* TG68K_ALU.vhd:379:24  */
  assign n9711 = exec[12]; // extract
  /* TG68K_ALU.vhd:380:47  */
  assign n9712 = bcd_pur[8]; // extract
  /* TG68K_ALU.vhd:380:36  */
  assign n9713 = ~n9712;
  /* TG68K_ALU.vhd:380:60  */
  assign n9714 = bcd_a[7]; // extract
  /* TG68K_ALU.vhd:380:51  */
  assign n9715 = n9713 & n9714;
  /* TG68K_ALU.vhd:382:41  */
  assign n9716 = bcd_pur[9:1]; // extract
  /* TG68K_ALU.vhd:382:54  */
  assign n9717 = n9716 + bcd_kor;
  /* TG68K_ALU.vhd:383:36  */
  assign n9718 = bcd_pur[4]; // extract
  /* TG68K_ALU.vhd:383:52  */
  assign n9719 = bcd_pur[3]; // extract
  /* TG68K_ALU.vhd:383:66  */
  assign n9720 = bcd_pur[2]; // extract
  /* TG68K_ALU.vhd:383:56  */
  assign n9721 = n9719 | n9720;
  /* TG68K_ALU.vhd:383:40  */
  assign n9722 = n9718 & n9721;
  /* TG68K_ALU.vhd:383:25  */
  assign n9724 = n9722 ? 4'b0110 : n9703;
  /* TG68K_ALU.vhd:386:36  */
  assign n9725 = bcd_pur[8]; // extract
  /* TG68K_ALU.vhd:386:52  */
  assign n9726 = bcd_pur[7]; // extract
  /* TG68K_ALU.vhd:386:66  */
  assign n9727 = bcd_pur[6]; // extract
  /* TG68K_ALU.vhd:386:56  */
  assign n9728 = n9726 | n9727;
  /* TG68K_ALU.vhd:386:81  */
  assign n9729 = bcd_pur[5]; // extract
  /* TG68K_ALU.vhd:386:96  */
  assign n9730 = bcd_pur[4]; // extract
  /* TG68K_ALU.vhd:386:85  */
  assign n9731 = n9729 & n9730;
  /* TG68K_ALU.vhd:386:112  */
  assign n9732 = bcd_pur[3]; // extract
  /* TG68K_ALU.vhd:386:126  */
  assign n9733 = bcd_pur[2]; // extract
  /* TG68K_ALU.vhd:386:116  */
  assign n9734 = n9732 | n9733;
  /* TG68K_ALU.vhd:386:100  */
  assign n9735 = n9731 & n9734;
  /* TG68K_ALU.vhd:386:70  */
  assign n9736 = n9728 | n9735;
  /* TG68K_ALU.vhd:386:40  */
  assign n9737 = n9725 & n9736;
  /* TG68K_ALU.vhd:386:25  */
  assign n9739 = n9737 ? 4'b0110 : n9709;
  /* TG68K_ALU.vhd:390:43  */
  assign n9740 = bcd_pur[8]; // extract
  /* TG68K_ALU.vhd:390:60  */
  assign n9741 = bcd_a[7]; // extract
  /* TG68K_ALU.vhd:390:51  */
  assign n9742 = ~n9741;
  /* TG68K_ALU.vhd:390:47  */
  assign n9743 = n9740 & n9742;
  /* TG68K_ALU.vhd:392:41  */
  assign n9744 = bcd_pur[9:1]; // extract
  /* TG68K_ALU.vhd:392:54  */
  assign n9745 = n9744 - bcd_kor;
  assign n9746 = {n9739, n9724};
  assign n9747 = {n9709, n9703};
  /* TG68K_ALU.vhd:379:17  */
  assign n9748 = n9711 ? n9746 : n9747;
  /* TG68K_ALU.vhd:379:17  */
  assign n9749 = n9711 ? n9715 : n9743;
  /* TG68K_ALU.vhd:379:17  */
  assign n9750 = n9711 ? n9717 : n9745;
  /* TG68K_ALU.vhd:394:23  */
  assign n9751 = cpu[1]; // extract
  /* TG68K_ALU.vhd:394:17  */
  assign n9753 = n9751 ? 1'b0 : n9749;
  /* TG68K_ALU.vhd:397:39  */
  assign n9754 = bcd_pur[9]; // extract
  /* TG68K_ALU.vhd:397:51  */
  assign n9755 = bcd_a[8]; // extract
  /* TG68K_ALU.vhd:397:43  */
  assign n9756 = n9754 | n9755;
  /* TG68K_ALU.vhd:409:44  */
  assign n9761 = opcode[7:6]; // extract
  /* TG68K_ALU.vhd:410:41  */
  assign n9763 = n9761 == 2'b01;
  /* TG68K_ALU.vhd:412:41  */
  assign n9765 = n9761 == 2'b11;
  assign n9766 = {n9765, n9763};
  /* TG68K_ALU.vhd:409:33  */
  always @*
    case (n9766)
      2'b10: n9769 = 1'b0;
      2'b01: n9769 = 1'b1;
      default: n9769 = 1'b0;
    endcase
  /* TG68K_ALU.vhd:409:33  */
  always @*
    case (n9766)
      2'b10: n9773 = 1'b1;
      2'b01: n9773 = 1'b0;
      default: n9773 = 1'b0;
    endcase
  /* TG68K_ALU.vhd:419:30  */
  assign n9779 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:419:33  */
  assign n9780 = ~n9779;
  /* TG68K_ALU.vhd:420:38  */
  assign n9781 = exe_opcode[5:4]; // extract
  /* TG68K_ALU.vhd:420:50  */
  assign n9783 = n9781 == 2'b00;
  /* TG68K_ALU.vhd:421:53  */
  assign n9784 = sndopc[4:0]; // extract
  /* TG68K_ALU.vhd:423:58  */
  assign n9785 = sndopc[2:0]; // extract
  /* TG68K_ALU.vhd:423:51  */
  assign n9787 = {2'b00, n9785};
  /* TG68K_ALU.vhd:420:25  */
  assign n9788 = n9783 ? n9784 : n9787;
  /* TG68K_ALU.vhd:426:38  */
  assign n9789 = exe_opcode[5:4]; // extract
  /* TG68K_ALU.vhd:426:50  */
  assign n9791 = n9789 == 2'b00;
  /* TG68K_ALU.vhd:427:53  */
  assign n9792 = reg_qb[4:0]; // extract
  /* TG68K_ALU.vhd:429:58  */
  assign n9793 = reg_qb[2:0]; // extract
  /* TG68K_ALU.vhd:429:51  */
  assign n9795 = {2'b00, n9793};
  /* TG68K_ALU.vhd:426:25  */
  assign n9796 = n9791 ? n9792 : n9795;
  /* TG68K_ALU.vhd:419:17  */
  assign n9797 = n9780 ? n9788 : n9796;
  /* TG68K_ALU.vhd:435:65  */
  assign n9803 = ~one_bit_in;
  /* TG68K_ALU.vhd:435:61  */
  assign n9804 = bchg & n9803;
  /* TG68K_ALU.vhd:435:81  */
  assign n9805 = n9804 | bset;
  /* TG68K_ALU.vhd:456:42  */
  assign n9811 = opcode[5:4]; // extract
  /* TG68K_ALU.vhd:456:55  */
  assign n9813 = n9811 == 2'b00;
  /* TG68K_ALU.vhd:456:33  */
  assign n9816 = n9813 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:459:44  */
  assign n9818 = opcode[10:8]; // extract
  /* TG68K_ALU.vhd:460:41  */
  assign n9820 = n9818 == 3'b010;
  /* TG68K_ALU.vhd:461:41  */
  assign n9822 = n9818 == 3'b011;
  /* TG68K_ALU.vhd:463:41  */
  assign n9824 = n9818 == 3'b101;
  /* TG68K_ALU.vhd:464:41  */
  assign n9826 = n9818 == 3'b110;
  /* TG68K_ALU.vhd:465:41  */
  assign n9828 = n9818 == 3'b111;
  assign n9829 = {n9828, n9826, n9824, n9822, n9820};
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n9829)
      5'b10000: n9832 = 1'b0;
      5'b01000: n9832 = 1'b1;
      5'b00100: n9832 = 1'b0;
      5'b00010: n9832 = 1'b0;
      5'b00001: n9832 = 1'b0;
      default: n9832 = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n9829)
      5'b10000: n9836 = 1'b0;
      5'b01000: n9836 = 1'b0;
      5'b00100: n9836 = 1'b0;
      5'b00010: n9836 = 1'b0;
      5'b00001: n9836 = 1'b1;
      default: n9836 = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n9829)
      5'b10000: n9840 = 1'b1;
      5'b01000: n9840 = 1'b0;
      5'b00100: n9840 = 1'b0;
      5'b00010: n9840 = 1'b0;
      5'b00001: n9840 = 1'b0;
      default: n9840 = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n9829)
      5'b10000: n9844 = 1'b0;
      5'b01000: n9844 = 1'b0;
      5'b00100: n9844 = 1'b0;
      5'b00010: n9844 = 1'b1;
      5'b00001: n9844 = 1'b0;
      default: n9844 = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n9829)
      5'b10000: n9848 = 1'b0;
      5'b01000: n9848 = 1'b0;
      5'b00100: n9848 = 1'b1;
      5'b00010: n9848 = 1'b0;
      5'b00001: n9848 = 1'b0;
      default: n9848 = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n9829)
      5'b10000: n9851 = 1'b1;
      5'b01000: n9851 = n9816;
      5'b00100: n9851 = n9816;
      5'b00010: n9851 = n9816;
      5'b00001: n9851 = n9816;
      default: n9851 = n9816;
    endcase
  /* TG68K_ALU.vhd:469:42  */
  assign n9852 = opcode[4:3]; // extract
  /* TG68K_ALU.vhd:469:54  */
  assign n9854 = n9852 == 2'b00;
  /* TG68K_ALU.vhd:469:33  */
  assign n9857 = n9854 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:472:53  */
  assign n9859 = result[39:32]; // extract
  /* TG68K_ALU.vhd:476:17  */
  assign n9876 = bf_ins ? reg_qb : bf_set2;
  /* TG68K_ALU.vhd:490:38  */
  assign n9877 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9879 = $unsigned(5'b00000) > $unsigned(n9877);
  assign n9882 = n9876[0]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9883 = n9879 ? 1'b0 : n9882;
  /* TG68K_ALU.vhd:490:25  */
  assign n9886 = n9879 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:490:38  */
  assign n9889 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9891 = $unsigned(5'b00001) > $unsigned(n9889);
  assign n9894 = n9876[1]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9895 = n9891 ? 1'b0 : n9894;
  assign n9897 = n9887[1]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9898 = n9891 ? 1'b1 : n9897;
  /* TG68K_ALU.vhd:490:38  */
  assign n9900 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9902 = $unsigned(5'b00010) > $unsigned(n9900);
  assign n9905 = n9876[2]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9906 = n9902 ? 1'b0 : n9905;
  assign n9908 = n9887[2]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9909 = n9902 ? 1'b1 : n9908;
  /* TG68K_ALU.vhd:490:38  */
  assign n9911 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9913 = $unsigned(5'b00011) > $unsigned(n9911);
  assign n9916 = n9876[3]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9917 = n9913 ? 1'b0 : n9916;
  assign n9919 = n9887[3]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9920 = n9913 ? 1'b1 : n9919;
  /* TG68K_ALU.vhd:490:38  */
  assign n9922 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9924 = $unsigned(5'b00100) > $unsigned(n9922);
  assign n9927 = n9876[4]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9928 = n9924 ? 1'b0 : n9927;
  assign n9930 = n9887[4]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9931 = n9924 ? 1'b1 : n9930;
  /* TG68K_ALU.vhd:490:38  */
  assign n9933 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9935 = $unsigned(5'b00101) > $unsigned(n9933);
  assign n9938 = n9876[5]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9939 = n9935 ? 1'b0 : n9938;
  assign n9941 = n9887[5]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9942 = n9935 ? 1'b1 : n9941;
  /* TG68K_ALU.vhd:490:38  */
  assign n9944 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9946 = $unsigned(5'b00110) > $unsigned(n9944);
  assign n9949 = n9876[6]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9950 = n9946 ? 1'b0 : n9949;
  assign n9952 = n9887[6]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9953 = n9946 ? 1'b1 : n9952;
  /* TG68K_ALU.vhd:490:38  */
  assign n9955 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9957 = $unsigned(5'b00111) > $unsigned(n9955);
  assign n9960 = n9876[7]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9961 = n9957 ? 1'b0 : n9960;
  assign n9963 = n9887[7]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9964 = n9957 ? 1'b1 : n9963;
  /* TG68K_ALU.vhd:490:38  */
  assign n9966 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9968 = $unsigned(5'b01000) > $unsigned(n9966);
  assign n9971 = n9876[8]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9972 = n9968 ? 1'b0 : n9971;
  assign n9974 = n9887[8]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9975 = n9968 ? 1'b1 : n9974;
  /* TG68K_ALU.vhd:490:38  */
  assign n9977 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9979 = $unsigned(5'b01001) > $unsigned(n9977);
  assign n9982 = n9876[9]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9983 = n9979 ? 1'b0 : n9982;
  assign n9985 = n9887[9]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9986 = n9979 ? 1'b1 : n9985;
  /* TG68K_ALU.vhd:490:38  */
  assign n9988 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n9990 = $unsigned(5'b01010) > $unsigned(n9988);
  assign n9993 = n9876[10]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9994 = n9990 ? 1'b0 : n9993;
  assign n9996 = n9887[10]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n9997 = n9990 ? 1'b1 : n9996;
  /* TG68K_ALU.vhd:490:38  */
  assign n9999 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10001 = $unsigned(5'b01011) > $unsigned(n9999);
  assign n10004 = n9876[11]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10005 = n10001 ? 1'b0 : n10004;
  assign n10007 = n9887[11]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10008 = n10001 ? 1'b1 : n10007;
  /* TG68K_ALU.vhd:490:38  */
  assign n10010 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10012 = $unsigned(5'b01100) > $unsigned(n10010);
  assign n10015 = n9876[12]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10016 = n10012 ? 1'b0 : n10015;
  assign n10018 = n9887[12]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10019 = n10012 ? 1'b1 : n10018;
  /* TG68K_ALU.vhd:490:38  */
  assign n10021 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10023 = $unsigned(5'b01101) > $unsigned(n10021);
  assign n10026 = n9876[13]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10027 = n10023 ? 1'b0 : n10026;
  assign n10029 = n9887[13]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10030 = n10023 ? 1'b1 : n10029;
  /* TG68K_ALU.vhd:490:38  */
  assign n10032 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10034 = $unsigned(5'b01110) > $unsigned(n10032);
  assign n10037 = n9876[14]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10038 = n10034 ? 1'b0 : n10037;
  assign n10040 = n9887[14]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10041 = n10034 ? 1'b1 : n10040;
  /* TG68K_ALU.vhd:490:38  */
  assign n10043 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10045 = $unsigned(5'b01111) > $unsigned(n10043);
  assign n10048 = n9876[15]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10049 = n10045 ? 1'b0 : n10048;
  assign n10051 = n9887[15]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10052 = n10045 ? 1'b1 : n10051;
  /* TG68K_ALU.vhd:490:38  */
  assign n10054 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10056 = $unsigned(5'b10000) > $unsigned(n10054);
  assign n10059 = n9876[16]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10060 = n10056 ? 1'b0 : n10059;
  assign n10062 = n9887[16]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10063 = n10056 ? 1'b1 : n10062;
  /* TG68K_ALU.vhd:490:38  */
  assign n10065 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10067 = $unsigned(5'b10001) > $unsigned(n10065);
  assign n10070 = n9876[17]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10071 = n10067 ? 1'b0 : n10070;
  assign n10073 = n9887[17]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10074 = n10067 ? 1'b1 : n10073;
  /* TG68K_ALU.vhd:490:38  */
  assign n10076 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10078 = $unsigned(5'b10010) > $unsigned(n10076);
  assign n10081 = n9876[18]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10082 = n10078 ? 1'b0 : n10081;
  assign n10084 = n9887[18]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10085 = n10078 ? 1'b1 : n10084;
  /* TG68K_ALU.vhd:490:38  */
  assign n10087 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10089 = $unsigned(5'b10011) > $unsigned(n10087);
  assign n10092 = n9876[19]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10093 = n10089 ? 1'b0 : n10092;
  assign n10095 = n9887[19]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10096 = n10089 ? 1'b1 : n10095;
  /* TG68K_ALU.vhd:490:38  */
  assign n10098 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10100 = $unsigned(5'b10100) > $unsigned(n10098);
  assign n10103 = n9876[20]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10104 = n10100 ? 1'b0 : n10103;
  assign n10106 = n9887[20]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10107 = n10100 ? 1'b1 : n10106;
  /* TG68K_ALU.vhd:490:38  */
  assign n10109 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10111 = $unsigned(5'b10101) > $unsigned(n10109);
  assign n10114 = n9876[21]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10115 = n10111 ? 1'b0 : n10114;
  assign n10117 = n9887[21]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10118 = n10111 ? 1'b1 : n10117;
  /* TG68K_ALU.vhd:490:38  */
  assign n10120 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10122 = $unsigned(5'b10110) > $unsigned(n10120);
  assign n10125 = n9876[22]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10126 = n10122 ? 1'b0 : n10125;
  assign n10128 = n9887[22]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10129 = n10122 ? 1'b1 : n10128;
  /* TG68K_ALU.vhd:490:38  */
  assign n10131 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10133 = $unsigned(5'b10111) > $unsigned(n10131);
  assign n10136 = n9876[23]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10137 = n10133 ? 1'b0 : n10136;
  assign n10139 = n9887[23]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10140 = n10133 ? 1'b1 : n10139;
  /* TG68K_ALU.vhd:490:38  */
  assign n10142 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10144 = $unsigned(5'b11000) > $unsigned(n10142);
  assign n10147 = n9876[24]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10148 = n10144 ? 1'b0 : n10147;
  assign n10150 = n9887[24]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10151 = n10144 ? 1'b1 : n10150;
  /* TG68K_ALU.vhd:490:38  */
  assign n10153 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10155 = $unsigned(5'b11001) > $unsigned(n10153);
  assign n10158 = n9876[25]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10159 = n10155 ? 1'b0 : n10158;
  assign n10161 = n9887[25]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10162 = n10155 ? 1'b1 : n10161;
  /* TG68K_ALU.vhd:490:38  */
  assign n10164 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10166 = $unsigned(5'b11010) > $unsigned(n10164);
  assign n10169 = n9876[26]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10170 = n10166 ? 1'b0 : n10169;
  assign n10172 = n9887[26]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10173 = n10166 ? 1'b1 : n10172;
  /* TG68K_ALU.vhd:490:38  */
  assign n10175 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10177 = $unsigned(5'b11011) > $unsigned(n10175);
  assign n10180 = n9876[27]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10181 = n10177 ? 1'b0 : n10180;
  assign n10183 = n9887[27]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10184 = n10177 ? 1'b1 : n10183;
  /* TG68K_ALU.vhd:490:38  */
  assign n10186 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10188 = $unsigned(5'b11100) > $unsigned(n10186);
  assign n10191 = n9876[28]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10192 = n10188 ? 1'b0 : n10191;
  assign n10194 = n9887[28]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10195 = n10188 ? 1'b1 : n10194;
  /* TG68K_ALU.vhd:490:38  */
  assign n10197 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10199 = $unsigned(5'b11101) > $unsigned(n10197);
  assign n10202 = n9876[29]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10203 = n10199 ? 1'b0 : n10202;
  assign n10205 = n9887[29]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10206 = n10199 ? 1'b1 : n10205;
  /* TG68K_ALU.vhd:490:38  */
  assign n10208 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10210 = $unsigned(5'b11110) > $unsigned(n10208);
  assign n10213 = n9876[30]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10214 = n10210 ? 1'b0 : n10213;
  assign n10215 = n9876[31]; // extract
  assign n10216 = n9887[30]; // extract
  /* TG68K_ALU.vhd:490:25  */
  assign n10217 = n10210 ? 1'b1 : n10216;
  assign n10218 = n9887[31]; // extract
  /* TG68K_ALU.vhd:490:38  */
  assign n10219 = bf_width[4:0]; // extract
  /* TG68K_ALU.vhd:490:29  */
  assign n10221 = $unsigned(5'b11111) > $unsigned(n10219);
  /* TG68K_ALU.vhd:490:25  */
  assign n10224 = n10221 ? 1'b0 : n10215;
  /* TG68K_ALU.vhd:490:25  */
  assign n10225 = n10221 ? 1'b1 : n10218;
  /* TG68K_ALU.vhd:496:37  */
  assign n10227 = bf_width[4:0];  // trunc
  /* TG68K_ALU.vhd:497:32  */
  assign n10230 = bf_nflag & bf_exts;
  /* TG68K_ALU.vhd:498:47  */
  assign n10231 = datareg | unshifted_bitmask;
  /* TG68K_ALU.vhd:497:17  */
  assign n10232 = n10230 ? n10231 : datareg;
  /* TG68K_ALU.vhd:504:30  */
  assign n10233 = bf_loffset[4]; // extract
  /* TG68K_ALU.vhd:505:57  */
  assign n10234 = unshifted_bitmask[15:0]; // extract
  /* TG68K_ALU.vhd:505:88  */
  assign n10235 = unshifted_bitmask[31:16]; // extract
  /* TG68K_ALU.vhd:505:70  */
  assign n10236 = {n10234, n10235};
  /* TG68K_ALU.vhd:504:17  */
  assign n10237 = n10233 ? n10236 : unshifted_bitmask;
  /* TG68K_ALU.vhd:509:30  */
  assign n10238 = bf_loffset[3]; // extract
  /* TG68K_ALU.vhd:510:64  */
  assign n10239 = bitmaskmux3[23:0]; // extract
  /* TG68K_ALU.vhd:510:89  */
  assign n10240 = bitmaskmux3[31:24]; // extract
  /* TG68K_ALU.vhd:510:77  */
  assign n10241 = {n10239, n10240};
  /* TG68K_ALU.vhd:509:17  */
  assign n10242 = n10238 ? n10241 : bitmaskmux3;
  /* TG68K_ALU.vhd:514:30  */
  assign n10243 = bf_loffset[2]; // extract
  /* TG68K_ALU.vhd:515:51  */
  assign n10245 = {bitmaskmux2, 4'b1111};
  /* TG68K_ALU.vhd:517:71  */
  assign n10246 = bitmaskmux2[31:28]; // extract
  assign n10247 = n10245[3:0]; // extract
  /* TG68K_ALU.vhd:516:25  */
  assign n10248 = bf_d32 ? n10246 : n10247;
  assign n10249 = n10245[35:4]; // extract
  /* TG68K_ALU.vhd:520:46  */
  assign n10251 = {4'b1111, bitmaskmux2};
  assign n10252 = {n10249, n10248};
  /* TG68K_ALU.vhd:514:17  */
  assign n10253 = n10243 ? n10252 : n10251;
  /* TG68K_ALU.vhd:522:30  */
  assign n10254 = bf_loffset[1]; // extract
  /* TG68K_ALU.vhd:523:51  */
  assign n10256 = {bitmaskmux1, 2'b11};
  /* TG68K_ALU.vhd:525:71  */
  assign n10257 = bitmaskmux1[31:30]; // extract
  assign n10258 = n10256[1:0]; // extract
  /* TG68K_ALU.vhd:524:25  */
  assign n10259 = bf_d32 ? n10257 : n10258;
  assign n10260 = n10256[37:2]; // extract
  /* TG68K_ALU.vhd:528:44  */
  assign n10262 = {2'b11, bitmaskmux1};
  assign n10263 = {n10260, n10259};
  /* TG68K_ALU.vhd:522:17  */
  assign n10264 = n10254 ? n10263 : n10262;
  /* TG68K_ALU.vhd:530:30  */
  assign n10265 = bf_loffset[0]; // extract
  /* TG68K_ALU.vhd:531:47  */
  assign n10267 = {1'b1, bitmaskmux0};
  /* TG68K_ALU.vhd:531:59  */
  assign n10269 = {n10267, 1'b1};
  /* TG68K_ALU.vhd:533:66  */
  assign n10270 = bitmaskmux0[31]; // extract
  assign n10271 = n10269[0]; // extract
  /* TG68K_ALU.vhd:532:25  */
  assign n10272 = bf_d32 ? n10270 : n10271;
  assign n10273 = n10269[39:1]; // extract
  /* TG68K_ALU.vhd:536:48  */
  assign n10275 = {2'b11, bitmaskmux0};
  assign n10276 = {n10273, n10272};
  /* TG68K_ALU.vhd:530:17  */
  assign n10277 = n10265 ? n10276 : n10275;
  /* TG68K_ALU.vhd:541:35  */
  assign n10278 = {bf_ext_in, op2out};
  /* TG68K_ALU.vhd:543:54  */
  assign n10279 = op2out[7:0]; // extract
  assign n10280 = n10278[39:32]; // extract
  /* TG68K_ALU.vhd:542:17  */
  assign n10281 = bf_s32 ? n10279 : n10280;
  assign n10282 = n10278[31:0]; // extract
  /* TG68K_ALU.vhd:546:28  */
  assign n10283 = bf_shift[0]; // extract
  /* TG68K_ALU.vhd:547:40  */
  assign n10284 = shift[0]; // extract
  /* TG68K_ALU.vhd:547:49  */
  assign n10285 = shift[39:1]; // extract
  /* TG68K_ALU.vhd:547:43  */
  assign n10286 = {n10284, n10285};
  /* TG68K_ALU.vhd:546:17  */
  assign n10287 = n10283 ? n10286 : shift;
  /* TG68K_ALU.vhd:551:28  */
  assign n10288 = bf_shift[1]; // extract
  /* TG68K_ALU.vhd:552:41  */
  assign n10289 = inmux0[1:0]; // extract
  /* TG68K_ALU.vhd:552:60  */
  assign n10290 = inmux0[39:2]; // extract
  /* TG68K_ALU.vhd:552:53  */
  assign n10291 = {n10289, n10290};
  /* TG68K_ALU.vhd:551:17  */
  assign n10292 = n10288 ? n10291 : inmux0;
  /* TG68K_ALU.vhd:556:28  */
  assign n10293 = bf_shift[2]; // extract
  /* TG68K_ALU.vhd:557:41  */
  assign n10294 = inmux1[3:0]; // extract
  /* TG68K_ALU.vhd:557:60  */
  assign n10295 = inmux1[39:4]; // extract
  /* TG68K_ALU.vhd:557:53  */
  assign n10296 = {n10294, n10295};
  /* TG68K_ALU.vhd:556:17  */
  assign n10297 = n10293 ? n10296 : inmux1;
  /* TG68K_ALU.vhd:561:28  */
  assign n10298 = bf_shift[3]; // extract
  /* TG68K_ALU.vhd:562:41  */
  assign n10299 = inmux2[7:0]; // extract
  /* TG68K_ALU.vhd:562:60  */
  assign n10300 = inmux2[31:8]; // extract
  /* TG68K_ALU.vhd:562:53  */
  assign n10301 = {n10299, n10300};
  /* TG68K_ALU.vhd:564:41  */
  assign n10302 = inmux2[31:0]; // extract
  /* TG68K_ALU.vhd:561:17  */
  assign n10303 = n10298 ? n10301 : n10302;
  /* TG68K_ALU.vhd:566:28  */
  assign n10304 = bf_shift[4]; // extract
  /* TG68K_ALU.vhd:567:55  */
  assign n10305 = inmux3[15:0]; // extract
  /* TG68K_ALU.vhd:567:75  */
  assign n10306 = inmux3[31:16]; // extract
  /* TG68K_ALU.vhd:567:68  */
  assign n10307 = {n10305, n10306};
  /* TG68K_ALU.vhd:566:17  */
  assign n10308 = n10304 ? n10307 : inmux3;
  /* TG68K_ALU.vhd:574:56  */
  assign n10309 = bf_set2[7:0]; // extract
  /* TG68K_ALU.vhd:576:48  */
  assign n10310 = ~op2out;
  /* TG68K_ALU.vhd:577:49  */
  assign n10311 = ~bf_ext_in;
  assign n10312 = {n10311, n10310};
  /* TG68K_ALU.vhd:575:17  */
  assign n10314 = bf_bchg ? n10312 : 40'b0000000000000000000000000000000000000000;
  assign n10315 = {n10309, bf_set2};
  /* TG68K_ALU.vhd:572:17  */
  assign n10316 = bf_ins ? n10315 : n10314;
  /* TG68K_ALU.vhd:581:17  */
  assign n10318 = bf_bset ? 40'b1111111111111111111111111111111111111111 : n10316;
  /* TG68K_ALU.vhd:586:48  */
  assign n10319 = {bf_ext_in, op1out};
  /* TG68K_ALU.vhd:588:48  */
  assign n10320 = {bf_ext_in, op2out};
  /* TG68K_ALU.vhd:585:17  */
  assign n10321 = bf_ins ? n10319 : n10320;
  /* TG68K_ALU.vhd:591:43  */
  assign n10322 = shifted_bitmask[0]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10323 = result_tmp[0]; // extract
  assign n10324 = n10318[0]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10325 = n10322 ? n10323 : n10324;
  /* TG68K_ALU.vhd:591:43  */
  assign n10327 = shifted_bitmask[1]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10328 = result_tmp[1]; // extract
  assign n10329 = n10318[1]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10330 = n10327 ? n10328 : n10329;
  /* TG68K_ALU.vhd:591:43  */
  assign n10332 = shifted_bitmask[2]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10333 = result_tmp[2]; // extract
  assign n10334 = n10318[2]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10335 = n10332 ? n10333 : n10334;
  /* TG68K_ALU.vhd:591:43  */
  assign n10337 = shifted_bitmask[3]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10338 = result_tmp[3]; // extract
  assign n10339 = n10318[3]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10340 = n10337 ? n10338 : n10339;
  /* TG68K_ALU.vhd:591:43  */
  assign n10342 = shifted_bitmask[4]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10343 = result_tmp[4]; // extract
  assign n10344 = n10318[4]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10345 = n10342 ? n10343 : n10344;
  /* TG68K_ALU.vhd:591:43  */
  assign n10347 = shifted_bitmask[5]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10348 = result_tmp[5]; // extract
  assign n10349 = n10318[5]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10350 = n10347 ? n10348 : n10349;
  /* TG68K_ALU.vhd:591:43  */
  assign n10352 = shifted_bitmask[6]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10353 = result_tmp[6]; // extract
  assign n10354 = n10318[6]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10355 = n10352 ? n10353 : n10354;
  /* TG68K_ALU.vhd:591:43  */
  assign n10357 = shifted_bitmask[7]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10358 = result_tmp[7]; // extract
  assign n10359 = n10318[7]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10360 = n10357 ? n10358 : n10359;
  /* TG68K_ALU.vhd:591:43  */
  assign n10362 = shifted_bitmask[8]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10363 = result_tmp[8]; // extract
  assign n10364 = n10318[8]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10365 = n10362 ? n10363 : n10364;
  /* TG68K_ALU.vhd:591:43  */
  assign n10367 = shifted_bitmask[9]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10368 = result_tmp[9]; // extract
  assign n10369 = n10318[9]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10370 = n10367 ? n10368 : n10369;
  /* TG68K_ALU.vhd:591:43  */
  assign n10372 = shifted_bitmask[10]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10373 = result_tmp[10]; // extract
  assign n10374 = n10318[10]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10375 = n10372 ? n10373 : n10374;
  /* TG68K_ALU.vhd:591:43  */
  assign n10377 = shifted_bitmask[11]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10378 = result_tmp[11]; // extract
  assign n10379 = n10318[11]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10380 = n10377 ? n10378 : n10379;
  /* TG68K_ALU.vhd:591:43  */
  assign n10382 = shifted_bitmask[12]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10383 = result_tmp[12]; // extract
  assign n10384 = n10318[12]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10385 = n10382 ? n10383 : n10384;
  /* TG68K_ALU.vhd:591:43  */
  assign n10387 = shifted_bitmask[13]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10388 = result_tmp[13]; // extract
  assign n10389 = n10318[13]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10390 = n10387 ? n10388 : n10389;
  /* TG68K_ALU.vhd:591:43  */
  assign n10392 = shifted_bitmask[14]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10393 = result_tmp[14]; // extract
  assign n10394 = n10318[14]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10395 = n10392 ? n10393 : n10394;
  /* TG68K_ALU.vhd:591:43  */
  assign n10397 = shifted_bitmask[15]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10398 = result_tmp[15]; // extract
  assign n10399 = n10318[15]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10400 = n10397 ? n10398 : n10399;
  /* TG68K_ALU.vhd:591:43  */
  assign n10402 = shifted_bitmask[16]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10403 = result_tmp[16]; // extract
  assign n10404 = n10318[16]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10405 = n10402 ? n10403 : n10404;
  /* TG68K_ALU.vhd:591:43  */
  assign n10407 = shifted_bitmask[17]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10408 = result_tmp[17]; // extract
  assign n10409 = n10318[17]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10410 = n10407 ? n10408 : n10409;
  /* TG68K_ALU.vhd:591:43  */
  assign n10412 = shifted_bitmask[18]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10413 = result_tmp[18]; // extract
  assign n10414 = n10318[18]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10415 = n10412 ? n10413 : n10414;
  /* TG68K_ALU.vhd:591:43  */
  assign n10417 = shifted_bitmask[19]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10418 = result_tmp[19]; // extract
  assign n10419 = n10318[19]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10420 = n10417 ? n10418 : n10419;
  /* TG68K_ALU.vhd:591:43  */
  assign n10422 = shifted_bitmask[20]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10423 = result_tmp[20]; // extract
  assign n10424 = n10318[20]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10425 = n10422 ? n10423 : n10424;
  /* TG68K_ALU.vhd:591:43  */
  assign n10427 = shifted_bitmask[21]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10428 = result_tmp[21]; // extract
  assign n10429 = n10318[21]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10430 = n10427 ? n10428 : n10429;
  /* TG68K_ALU.vhd:591:43  */
  assign n10432 = shifted_bitmask[22]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10433 = result_tmp[22]; // extract
  assign n10434 = n10318[22]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10435 = n10432 ? n10433 : n10434;
  /* TG68K_ALU.vhd:591:43  */
  assign n10437 = shifted_bitmask[23]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10438 = result_tmp[23]; // extract
  assign n10439 = n10318[23]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10440 = n10437 ? n10438 : n10439;
  /* TG68K_ALU.vhd:591:43  */
  assign n10442 = shifted_bitmask[24]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10443 = result_tmp[24]; // extract
  assign n10444 = n10318[24]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10445 = n10442 ? n10443 : n10444;
  /* TG68K_ALU.vhd:591:43  */
  assign n10447 = shifted_bitmask[25]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10448 = result_tmp[25]; // extract
  assign n10449 = n10318[25]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10450 = n10447 ? n10448 : n10449;
  /* TG68K_ALU.vhd:591:43  */
  assign n10452 = shifted_bitmask[26]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10453 = result_tmp[26]; // extract
  assign n10454 = n10318[26]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10455 = n10452 ? n10453 : n10454;
  /* TG68K_ALU.vhd:591:43  */
  assign n10457 = shifted_bitmask[27]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10458 = result_tmp[27]; // extract
  assign n10459 = n10318[27]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10460 = n10457 ? n10458 : n10459;
  /* TG68K_ALU.vhd:591:43  */
  assign n10462 = shifted_bitmask[28]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10463 = result_tmp[28]; // extract
  assign n10464 = n10318[28]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10465 = n10462 ? n10463 : n10464;
  /* TG68K_ALU.vhd:591:43  */
  assign n10467 = shifted_bitmask[29]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10468 = result_tmp[29]; // extract
  assign n10469 = n10318[29]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10470 = n10467 ? n10468 : n10469;
  /* TG68K_ALU.vhd:591:43  */
  assign n10472 = shifted_bitmask[30]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10473 = result_tmp[30]; // extract
  assign n10474 = n10318[30]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10475 = n10472 ? n10473 : n10474;
  /* TG68K_ALU.vhd:591:43  */
  assign n10477 = shifted_bitmask[31]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10478 = result_tmp[31]; // extract
  assign n10479 = n10318[31]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10480 = n10477 ? n10478 : n10479;
  /* TG68K_ALU.vhd:591:43  */
  assign n10482 = shifted_bitmask[32]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10483 = result_tmp[32]; // extract
  assign n10484 = n10318[32]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10485 = n10482 ? n10483 : n10484;
  /* TG68K_ALU.vhd:591:43  */
  assign n10487 = shifted_bitmask[33]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10488 = result_tmp[33]; // extract
  assign n10489 = n10318[33]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10490 = n10487 ? n10488 : n10489;
  /* TG68K_ALU.vhd:591:43  */
  assign n10492 = shifted_bitmask[34]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10493 = result_tmp[34]; // extract
  assign n10494 = n10318[34]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10495 = n10492 ? n10493 : n10494;
  /* TG68K_ALU.vhd:591:43  */
  assign n10497 = shifted_bitmask[35]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10498 = result_tmp[35]; // extract
  assign n10499 = n10318[35]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10500 = n10497 ? n10498 : n10499;
  /* TG68K_ALU.vhd:591:43  */
  assign n10502 = shifted_bitmask[36]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10503 = result_tmp[36]; // extract
  assign n10504 = n10318[36]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10505 = n10502 ? n10503 : n10504;
  /* TG68K_ALU.vhd:591:43  */
  assign n10507 = shifted_bitmask[37]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10508 = result_tmp[37]; // extract
  assign n10509 = n10318[37]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10510 = n10507 ? n10508 : n10509;
  /* TG68K_ALU.vhd:591:43  */
  assign n10512 = shifted_bitmask[38]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10513 = result_tmp[38]; // extract
  assign n10514 = n10318[38]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10515 = n10512 ? n10513 : n10514;
  assign n10516 = n10318[39]; // extract
  /* TG68K_ALU.vhd:591:43  */
  assign n10517 = shifted_bitmask[39]; // extract
  /* TG68K_ALU.vhd:592:56  */
  assign n10518 = result_tmp[39]; // extract
  /* TG68K_ALU.vhd:591:25  */
  assign n10519 = n10517 ? n10518 : n10516;
  /* TG68K_ALU.vhd:598:36  */
  assign n10521 = {1'b0, bitnr};
  /* TG68K_ALU.vhd:598:43  */
  assign n10522 = {5'b0, mask_not_zero};  //  uext
  /* TG68K_ALU.vhd:598:43  */
  assign n10523 = n10521 + n10522;
  /* TG68K_ALU.vhd:601:24  */
  assign n10524 = mask[31:28]; // extract
  /* TG68K_ALU.vhd:601:38  */
  assign n10526 = n10524 == 4'b0000;
  /* TG68K_ALU.vhd:602:32  */
  assign n10527 = mask[27:24]; // extract
  /* TG68K_ALU.vhd:602:46  */
  assign n10529 = n10527 == 4'b0000;
  /* TG68K_ALU.vhd:603:40  */
  assign n10530 = mask[23:20]; // extract
  /* TG68K_ALU.vhd:603:54  */
  assign n10532 = n10530 == 4'b0000;
  /* TG68K_ALU.vhd:604:48  */
  assign n10533 = mask[19:16]; // extract
  /* TG68K_ALU.vhd:604:62  */
  assign n10535 = n10533 == 4'b0000;
  /* TG68K_ALU.vhd:606:56  */
  assign n10537 = mask[15:12]; // extract
  /* TG68K_ALU.vhd:606:70  */
  assign n10539 = n10537 == 4'b0000;
  /* TG68K_ALU.vhd:607:64  */
  assign n10540 = mask[11:8]; // extract
  /* TG68K_ALU.vhd:607:77  */
  assign n10542 = n10540 == 4'b0000;
  /* TG68K_ALU.vhd:609:72  */
  assign n10544 = mask[7:4]; // extract
  /* TG68K_ALU.vhd:609:84  */
  assign n10546 = n10544 == 4'b0000;
  /* TG68K_ALU.vhd:611:84  */
  assign n10548 = mask[3:0]; // extract
  /* TG68K_ALU.vhd:613:84  */
  assign n10549 = mask[7:4]; // extract
  /* TG68K_ALU.vhd:609:65  */
  assign n10550 = n10546 ? n10548 : n10549;
  /* TG68K_ALU.vhd:609:65  */
  assign n10552 = n10546 ? 1'b0 : 1'b1;
  /* TG68K_ALU.vhd:616:76  */
  assign n10553 = mask[11:8]; // extract
  /* TG68K_ALU.vhd:607:57  */
  assign n10555 = n10542 ? n10550 : n10553;
  assign n10556 = {1'b0, n10552};
  assign n10557 = n10556[0]; // extract
  /* TG68K_ALU.vhd:607:57  */
  assign n10558 = n10542 ? n10557 : 1'b0;
  assign n10559 = n10556[1]; // extract
  /* TG68K_ALU.vhd:607:57  */
  assign n10561 = n10542 ? n10559 : 1'b1;
  /* TG68K_ALU.vhd:620:68  */
  assign n10562 = mask[15:12]; // extract
  /* TG68K_ALU.vhd:606:49  */
  assign n10563 = n10539 ? n10555 : n10562;
  assign n10564 = {n10561, n10558};
  /* TG68K_ALU.vhd:606:49  */
  assign n10566 = n10539 ? n10564 : 2'b11;
  /* TG68K_ALU.vhd:623:60  */
  assign n10567 = mask[19:16]; // extract
  /* TG68K_ALU.vhd:604:41  */
  assign n10570 = n10535 ? n10563 : n10567;
  assign n10571 = {1'b0, 1'b0};
  assign n10572 = {1'b0, n10566};
  assign n10573 = n10572[1:0]; // extract
  /* TG68K_ALU.vhd:604:41  */
  assign n10574 = n10535 ? n10573 : n10571;
  assign n10575 = n10572[2]; // extract
  /* TG68K_ALU.vhd:604:41  */
  assign n10577 = n10535 ? n10575 : 1'b1;
  /* TG68K_ALU.vhd:628:52  */
  assign n10578 = mask[23:20]; // extract
  /* TG68K_ALU.vhd:603:33  */
  assign n10580 = n10532 ? n10570 : n10578;
  assign n10581 = {n10577, n10574};
  assign n10582 = n10581[0]; // extract
  /* TG68K_ALU.vhd:603:33  */
  assign n10584 = n10532 ? n10582 : 1'b1;
  assign n10585 = n10581[1]; // extract
  /* TG68K_ALU.vhd:603:33  */
  assign n10586 = n10532 ? n10585 : 1'b0;
  assign n10587 = n10581[2]; // extract
  /* TG68K_ALU.vhd:603:33  */
  assign n10589 = n10532 ? n10587 : 1'b1;
  /* TG68K_ALU.vhd:632:44  */
  assign n10590 = mask[27:24]; // extract
  /* TG68K_ALU.vhd:602:25  */
  assign n10592 = n10529 ? n10580 : n10590;
  assign n10593 = {n10589, n10586, n10584};
  assign n10594 = n10593[0]; // extract
  /* TG68K_ALU.vhd:602:25  */
  assign n10595 = n10529 ? n10594 : 1'b0;
  assign n10596 = n10593[2:1]; // extract
  /* TG68K_ALU.vhd:602:25  */
  assign n10598 = n10529 ? n10596 : 2'b11;
  /* TG68K_ALU.vhd:636:36  */
  assign n10599 = mask[31:28]; // extract
  /* TG68K_ALU.vhd:601:17  */
  assign n10600 = n10526 ? n10592 : n10599;
  assign n10601 = {n10598, n10595};
  /* TG68K_ALU.vhd:601:17  */
  assign n10603 = n10526 ? n10601 : 3'b111;
  /* TG68K_ALU.vhd:639:23  */
  assign n10606 = mux[3:2]; // extract
  /* TG68K_ALU.vhd:639:35  */
  assign n10608 = n10606 == 2'b00;
  /* TG68K_ALU.vhd:641:31  */
  assign n10610 = mux[1]; // extract
  /* TG68K_ALU.vhd:641:34  */
  assign n10611 = ~n10610;
  /* TG68K_ALU.vhd:643:39  */
  assign n10613 = mux[0]; // extract
  /* TG68K_ALU.vhd:643:42  */
  assign n10614 = ~n10613;
  /* TG68K_ALU.vhd:643:33  */
  assign n10617 = n10614 ? 1'b0 : 1'b1;
  assign n10618 = n10604[0]; // extract
  /* TG68K_ALU.vhd:641:25  */
  assign n10619 = n10611 ? 1'b0 : n10618;
  /* TG68K_ALU.vhd:641:25  */
  assign n10621 = n10611 ? n10617 : 1'b1;
  /* TG68K_ALU.vhd:648:31  */
  assign n10622 = mux[3]; // extract
  /* TG68K_ALU.vhd:648:34  */
  assign n10623 = ~n10622;
  assign n10625 = n10604[0]; // extract
  /* TG68K_ALU.vhd:648:25  */
  assign n10626 = n10623 ? 1'b0 : n10625;
  assign n10627 = {1'b0, n10619};
  assign n10628 = n10627[0]; // extract
  /* TG68K_ALU.vhd:639:17  */
  assign n10629 = n10608 ? n10628 : n10626;
  assign n10630 = n10627[1]; // extract
  assign n10631 = n10604[1]; // extract
  /* TG68K_ALU.vhd:639:17  */
  assign n10632 = n10608 ? n10630 : n10631;
  /* TG68K_ALU.vhd:639:17  */
  assign n10635 = n10608 ? n10621 : 1'b1;
  /* TG68K_ALU.vhd:659:32  */
  assign n10640 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:661:66  */
  assign n10641 = op1out[7]; // extract
  /* TG68K_ALU.vhd:660:25  */
  assign n10643 = n10640 == 2'b00;
  /* TG68K_ALU.vhd:663:66  */
  assign n10644 = op1out[15]; // extract
  /* TG68K_ALU.vhd:662:25  */
  assign n10646 = n10640 == 2'b01;
  /* TG68K_ALU.vhd:662:34  */
  assign n10648 = n10640 == 2'b11;
  /* TG68K_ALU.vhd:662:34  */
  assign n10649 = n10646 | n10648;
  /* TG68K_ALU.vhd:665:66  */
  assign n10650 = op1out[31]; // extract
  /* TG68K_ALU.vhd:664:25  */
  assign n10652 = n10640 == 2'b10;
  assign n10653 = {n10652, n10649, n10643};
  /* TG68K_ALU.vhd:659:17  */
  always @*
    case (n10653)
      3'b100: n10654 = n10650;
      3'b010: n10654 = n10644;
      3'b001: n10654 = n10641;
      default: n10654 = rot_rot;
    endcase
  /* TG68K_ALU.vhd:685:24  */
  assign n10672 = exec[23]; // extract
  /* TG68K_ALU.vhd:687:39  */
  assign n10673 = n11806[4]; // extract
  /* TG68K_ALU.vhd:688:36  */
  assign n10675 = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:689:47  */
  assign n10676 = n11806[4]; // extract
  /* TG68K_ALU.vhd:688:25  */
  assign n10678 = n10675 ? n10676 : 1'b0;
  /* TG68K_ALU.vhd:694:38  */
  assign n10679 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:699:48  */
  assign n10682 = op1out[0]; // extract
  /* TG68K_ALU.vhd:700:48  */
  assign n10683 = op1out[0]; // extract
  /* TG68K_ALU.vhd:694:25  */
  assign n10703 = n10679 ? rot_rot : n10682;
  /* TG68K_ALU.vhd:694:25  */
  assign n10704 = n10679 ? rot_rot : n10683;
  /* TG68K_ALU.vhd:685:17  */
  assign n10707 = n10672 ? n10673 : n10703;
  /* TG68K_ALU.vhd:685:17  */
  assign n10708 = n10672 ? n10678 : n10704;
  /* TG68K_ALU.vhd:685:17  */
  assign n10709 = n10672 ? op1out : bsout;
  /* TG68K_ALU.vhd:723:28  */
  assign n10714 = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:724:40  */
  assign n10715 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:725:33  */
  assign n10717 = n10715 == 2'b00;
  /* TG68K_ALU.vhd:727:33  */
  assign n10719 = n10715 == 2'b01;
  /* TG68K_ALU.vhd:727:42  */
  assign n10721 = n10715 == 2'b11;
  /* TG68K_ALU.vhd:727:42  */
  assign n10722 = n10719 | n10721;
  /* TG68K_ALU.vhd:729:33  */
  assign n10724 = n10715 == 2'b10;
  assign n10725 = {n10724, n10722, n10717};
  /* TG68K_ALU.vhd:724:25  */
  always @*
    case (n10725)
      3'b100: n10730 = 6'b100001;
      3'b010: n10730 = 6'b010001;
      3'b001: n10730 = 6'b001001;
      default: n10730 = 6'b100000;
    endcase
  /* TG68K_ALU.vhd:734:40  */
  assign n10731 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:735:33  */
  assign n10733 = n10731 == 2'b00;
  /* TG68K_ALU.vhd:737:33  */
  assign n10735 = n10731 == 2'b01;
  /* TG68K_ALU.vhd:737:42  */
  assign n10737 = n10731 == 2'b11;
  /* TG68K_ALU.vhd:737:42  */
  assign n10738 = n10735 | n10737;
  /* TG68K_ALU.vhd:739:33  */
  assign n10740 = n10731 == 2'b10;
  assign n10741 = {n10740, n10738, n10733};
  /* TG68K_ALU.vhd:734:25  */
  always @*
    case (n10741)
      3'b100: n10746 = 6'b100000;
      3'b010: n10746 = 6'b010000;
      3'b001: n10746 = 6'b001000;
      default: n10746 = 6'b100000;
    endcase
  /* TG68K_ALU.vhd:723:17  */
  assign n10747 = n10714 ? n10730 : n10746;
  /* TG68K_ALU.vhd:745:30  */
  assign n10749 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:745:42  */
  assign n10751 = n10749 == 2'b11;
  /* TG68K_ALU.vhd:745:55  */
  assign n10752 = exec[81]; // extract
  /* TG68K_ALU.vhd:745:64  */
  assign n10753 = ~n10752;
  /* TG68K_ALU.vhd:745:48  */
  assign n10754 = n10751 | n10753;
  /* TG68K_ALU.vhd:747:33  */
  assign n10755 = exe_opcode[5]; // extract
  /* TG68K_ALU.vhd:748:43  */
  assign n10756 = op2out[5:0]; // extract
  /* TG68K_ALU.vhd:750:59  */
  assign n10757 = exe_opcode[11:9]; // extract
  /* TG68K_ALU.vhd:751:38  */
  assign n10758 = exe_opcode[11:9]; // extract
  /* TG68K_ALU.vhd:751:51  */
  assign n10760 = n10758 == 3'b000;
  /* TG68K_ALU.vhd:751:25  */
  assign n10763 = n10760 ? 3'b001 : 3'b000;
  assign n10764 = {n10763, n10757};
  /* TG68K_ALU.vhd:747:17  */
  assign n10765 = n10755 ? n10756 : n10764;
  /* TG68K_ALU.vhd:745:17  */
  assign n10767 = n10754 ? 6'b000001 : n10765;
  /* TG68K_ALU.vhd:762:29  */
  assign n10774 = $unsigned(bs_shift) < $unsigned(ring);
  /* TG68K_ALU.vhd:763:40  */
  assign n10775 = ring - bs_shift;
  /* TG68K_ALU.vhd:762:17  */
  assign n10777 = n10774 ? n10775 : 6'b000000;
  /* TG68K_ALU.vhd:765:45  */
  assign n10779 = vector[30:0]; // extract
  /* TG68K_ALU.vhd:765:38  */
  assign n10781 = {1'b0, n10779};
  /* TG68K_ALU.vhd:765:75  */
  assign n10782 = vector[31:1]; // extract
  /* TG68K_ALU.vhd:765:68  */
  assign n10784 = {1'b0, n10782};
  /* TG68K_ALU.vhd:765:60  */
  assign n10785 = n10781 ^ n10784;
  /* TG68K_ALU.vhd:765:90  */
  assign n10786 = {n10785, msb};
  /* TG68K_ALU.vhd:766:32  */
  assign n10787 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:767:25  */
  assign n10790 = n10787 == 2'b00;
  /* TG68K_ALU.vhd:769:25  */
  assign n10793 = n10787 == 2'b01;
  /* TG68K_ALU.vhd:769:34  */
  assign n10795 = n10787 == 2'b11;
  /* TG68K_ALU.vhd:769:34  */
  assign n10796 = n10793 | n10795;
  assign n10797 = {n10796, n10790};
  assign n10798 = n10786[8]; // extract
  /* TG68K_ALU.vhd:766:17  */
  always @*
    case (n10797)
      2'b10: n10799 = n10798;
      2'b01: n10799 = 1'b0;
      default: n10799 = n10798;
    endcase
  assign n10800 = n10786[16]; // extract
  /* TG68K_ALU.vhd:766:17  */
  always @*
    case (n10797)
      2'b10: n10801 = 1'b0;
      2'b01: n10801 = n10800;
      default: n10801 = n10800;
    endcase
  assign n10803 = n10786[7:0]; // extract
  assign n10804 = n10786[32:17]; // extract
  assign n10805 = n10786[15:9]; // extract
  /* TG68K_ALU.vhd:773:56  */
  assign n10806 = hot_msb[31:0]; // extract
  /* TG68K_ALU.vhd:773:48  */
  assign n10808 = {1'b0, n10806};
  /* TG68K_ALU.vhd:773:42  */
  assign n10809 = asl_over_xor - n10808;
  /* TG68K_ALU.vhd:775:28  */
  assign n10811 = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:775:48  */
  assign n10812 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:775:34  */
  assign n10813 = n10812 & n10811;
  /* TG68K_ALU.vhd:776:45  */
  assign n10814 = asl_over[32]; // extract
  /* TG68K_ALU.vhd:776:33  */
  assign n10815 = ~n10814;
  /* TG68K_ALU.vhd:775:17  */
  assign n10817 = n10813 ? n10815 : 1'b0;
  /* TG68K_ALU.vhd:780:30  */
  assign n10819 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:780:33  */
  assign n10820 = ~n10819;
  /* TG68K_ALU.vhd:781:42  */
  assign n10821 = result_bs[31]; // extract
  /* TG68K_ALU.vhd:783:40  */
  assign n10822 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:785:58  */
  assign n10823 = result_bs[8]; // extract
  /* TG68K_ALU.vhd:784:33  */
  assign n10825 = n10822 == 2'b00;
  /* TG68K_ALU.vhd:787:58  */
  assign n10826 = result_bs[16]; // extract
  /* TG68K_ALU.vhd:786:33  */
  assign n10828 = n10822 == 2'b01;
  /* TG68K_ALU.vhd:786:42  */
  assign n10830 = n10822 == 2'b11;
  /* TG68K_ALU.vhd:786:42  */
  assign n10831 = n10828 | n10830;
  /* TG68K_ALU.vhd:789:58  */
  assign n10832 = result_bs[32]; // extract
  /* TG68K_ALU.vhd:788:33  */
  assign n10834 = n10822 == 2'b10;
  assign n10835 = {n10834, n10831, n10825};
  /* TG68K_ALU.vhd:783:25  */
  always @*
    case (n10835)
      3'b100: n10836 = n10832;
      3'b010: n10836 = n10826;
      3'b001: n10836 = n10823;
      default: n10836 = bs_c;
    endcase
  /* TG68K_ALU.vhd:780:17  */
  assign n10837 = n10820 ? n10821 : n10836;
  /* TG68K_ALU.vhd:795:28  */
  assign n10839 = rot_bits == 2'b11;
  /* TG68K_ALU.vhd:796:38  */
  assign n10840 = n11806[4]; // extract
  /* TG68K_ALU.vhd:797:40  */
  assign n10841 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:799:69  */
  assign n10842 = result_bs[7:0]; // extract
  /* TG68K_ALU.vhd:799:94  */
  assign n10843 = result_bs[15:8]; // extract
  /* TG68K_ALU.vhd:799:82  */
  assign n10844 = n10842 | n10843;
  /* TG68K_ALU.vhd:800:52  */
  assign n10845 = alu[7]; // extract
  /* TG68K_ALU.vhd:798:33  */
  assign n10847 = n10841 == 2'b00;
  /* TG68K_ALU.vhd:802:70  */
  assign n10848 = result_bs[15:0]; // extract
  /* TG68K_ALU.vhd:802:96  */
  assign n10849 = result_bs[31:16]; // extract
  /* TG68K_ALU.vhd:802:84  */
  assign n10850 = n10848 | n10849;
  /* TG68K_ALU.vhd:803:52  */
  assign n10851 = alu[15]; // extract
  /* TG68K_ALU.vhd:801:33  */
  assign n10853 = n10841 == 2'b01;
  /* TG68K_ALU.vhd:801:42  */
  assign n10855 = n10841 == 2'b11;
  /* TG68K_ALU.vhd:801:42  */
  assign n10856 = n10853 | n10855;
  /* TG68K_ALU.vhd:805:57  */
  assign n10857 = result_bs[31:0]; // extract
  /* TG68K_ALU.vhd:805:83  */
  assign n10858 = result_bs[63:32]; // extract
  /* TG68K_ALU.vhd:805:71  */
  assign n10859 = n10857 | n10858;
  /* TG68K_ALU.vhd:806:52  */
  assign n10860 = alu[31]; // extract
  /* TG68K_ALU.vhd:804:33  */
  assign n10862 = n10841 == 2'b10;
  assign n10863 = {n10862, n10856, n10847};
  assign n10864 = n10850[7:0]; // extract
  assign n10865 = n10859[7:0]; // extract
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n10863)
      3'b100: n10867 = n10865;
      3'b010: n10867 = n10864;
      3'b001: n10867 = n10844;
      default: n10867 = 8'bX;
    endcase
  assign n10868 = n10850[15:8]; // extract
  assign n10869 = n10859[15:8]; // extract
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n10863)
      3'b100: n10871 = n10869;
      3'b010: n10871 = n10868;
      3'b001: n10871 = 8'bX;
      default: n10871 = 8'bX;
    endcase
  assign n10872 = n10859[31:16]; // extract
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n10863)
      3'b100: n10874 = n10872;
      3'b010: n10874 = 16'bX;
      3'b001: n10874 = 16'bX;
      default: n10874 = 16'bX;
    endcase
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n10863)
      3'b100: n10875 = n10860;
      3'b010: n10875 = n10851;
      3'b001: n10875 = n10845;
      default: n10875 = n10837;
    endcase
  /* TG68K_ALU.vhd:809:38  */
  assign n10876 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:810:44  */
  assign n10877 = alu[0]; // extract
  /* TG68K_ALU.vhd:809:25  */
  assign n10878 = n10876 ? n10877 : n10875;
  /* TG68K_ALU.vhd:812:31  */
  assign n10880 = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:813:40  */
  assign n10881 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:815:69  */
  assign n10882 = result_bs[7:0]; // extract
  /* TG68K_ALU.vhd:815:94  */
  assign n10883 = result_bs[16:9]; // extract
  /* TG68K_ALU.vhd:815:82  */
  assign n10884 = n10882 | n10883;
  /* TG68K_ALU.vhd:816:58  */
  assign n10885 = result_bs[8]; // extract
  /* TG68K_ALU.vhd:816:74  */
  assign n10886 = result_bs[17]; // extract
  /* TG68K_ALU.vhd:816:62  */
  assign n10887 = n10885 | n10886;
  /* TG68K_ALU.vhd:814:33  */
  assign n10889 = n10881 == 2'b00;
  /* TG68K_ALU.vhd:818:70  */
  assign n10890 = result_bs[15:0]; // extract
  /* TG68K_ALU.vhd:818:96  */
  assign n10891 = result_bs[32:17]; // extract
  /* TG68K_ALU.vhd:818:84  */
  assign n10892 = n10890 | n10891;
  /* TG68K_ALU.vhd:819:58  */
  assign n10893 = result_bs[16]; // extract
  /* TG68K_ALU.vhd:819:75  */
  assign n10894 = result_bs[33]; // extract
  /* TG68K_ALU.vhd:819:63  */
  assign n10895 = n10893 | n10894;
  /* TG68K_ALU.vhd:817:33  */
  assign n10897 = n10881 == 2'b01;
  /* TG68K_ALU.vhd:817:42  */
  assign n10899 = n10881 == 2'b11;
  /* TG68K_ALU.vhd:817:42  */
  assign n10900 = n10897 | n10899;
  /* TG68K_ALU.vhd:821:57  */
  assign n10901 = result_bs[31:0]; // extract
  /* TG68K_ALU.vhd:821:83  */
  assign n10902 = result_bs[64:33]; // extract
  /* TG68K_ALU.vhd:821:71  */
  assign n10903 = n10901 | n10902;
  /* TG68K_ALU.vhd:822:58  */
  assign n10904 = result_bs[32]; // extract
  /* TG68K_ALU.vhd:822:75  */
  assign n10905 = result_bs[65]; // extract
  /* TG68K_ALU.vhd:822:63  */
  assign n10906 = n10904 | n10905;
  /* TG68K_ALU.vhd:820:33  */
  assign n10908 = n10881 == 2'b10;
  assign n10909 = {n10908, n10900, n10889};
  assign n10910 = n10892[7:0]; // extract
  assign n10911 = n10903[7:0]; // extract
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n10909)
      3'b100: n10913 = n10911;
      3'b010: n10913 = n10910;
      3'b001: n10913 = n10884;
      default: n10913 = 8'bX;
    endcase
  assign n10914 = n10892[15:8]; // extract
  assign n10915 = n10903[15:8]; // extract
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n10909)
      3'b100: n10917 = n10915;
      3'b010: n10917 = n10914;
      3'b001: n10917 = 8'bX;
      default: n10917 = 8'bX;
    endcase
  assign n10918 = n10903[31:16]; // extract
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n10909)
      3'b100: n10920 = n10918;
      3'b010: n10920 = 16'bX;
      3'b001: n10920 = 16'bX;
      default: n10920 = 16'bX;
    endcase
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n10909)
      3'b100: n10921 = n10906;
      3'b010: n10921 = n10895;
      3'b001: n10921 = n10887;
      default: n10921 = n10837;
    endcase
  /* TG68K_ALU.vhd:826:38  */
  assign n10922 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:826:41  */
  assign n10923 = ~n10922;
  /* TG68K_ALU.vhd:827:49  */
  assign n10924 = result_bs[63:32]; // extract
  /* TG68K_ALU.vhd:829:49  */
  assign n10925 = result_bs[31:0]; // extract
  /* TG68K_ALU.vhd:826:25  */
  assign n10926 = n10923 ? n10924 : n10925;
  assign n10927 = {n10920, n10917, n10913};
  /* TG68K_ALU.vhd:812:17  */
  assign n10928 = n10880 ? n10927 : n10926;
  /* TG68K_ALU.vhd:812:17  */
  assign n10929 = n10880 ? n10921 : n10837;
  assign n10930 = {n10874, n10871, n10867};
  /* TG68K_ALU.vhd:795:17  */
  assign n10931 = n10839 ? n10930 : n10928;
  /* TG68K_ALU.vhd:795:17  */
  assign n10933 = n10839 ? n10878 : n10929;
  /* TG68K_ALU.vhd:795:17  */
  assign n10934 = n10839 ? n10840 : bs_c;
  /* TG68K_ALU.vhd:833:29  */
  assign n10936 = bs_shift == 6'b000000;
  /* TG68K_ALU.vhd:834:36  */
  assign n10938 = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:835:46  */
  assign n10939 = n11806[4]; // extract
  /* TG68K_ALU.vhd:834:25  */
  assign n10941 = n10938 ? n10939 : 1'b0;
  /* TG68K_ALU.vhd:839:38  */
  assign n10942 = n11806[4]; // extract
  /* TG68K_ALU.vhd:833:17  */
  assign n10944 = n10936 ? 1'b0 : n10817;
  /* TG68K_ALU.vhd:833:17  */
  assign n10945 = n10936 ? n10941 : n10933;
  /* TG68K_ALU.vhd:833:17  */
  assign n10946 = n10936 ? n10942 : n10934;
  /* TG68K_ALU.vhd:848:45  */
  assign n10948 = bs_shift == 6'b111111;
  /* TG68K_ALU.vhd:850:48  */
  assign n10950 = $unsigned(bs_shift) > $unsigned(6'b110101);
  /* TG68K_ALU.vhd:851:66  */
  assign n10952 = bs_shift - 6'b110110;
  /* TG68K_ALU.vhd:852:48  */
  assign n10954 = $unsigned(bs_shift) > $unsigned(6'b101100);
  /* TG68K_ALU.vhd:853:66  */
  assign n10956 = bs_shift - 6'b101101;
  /* TG68K_ALU.vhd:854:48  */
  assign n10958 = $unsigned(bs_shift) > $unsigned(6'b100011);
  /* TG68K_ALU.vhd:855:66  */
  assign n10960 = bs_shift - 6'b100100;
  /* TG68K_ALU.vhd:856:48  */
  assign n10962 = $unsigned(bs_shift) > $unsigned(6'b011010);
  /* TG68K_ALU.vhd:857:66  */
  assign n10964 = bs_shift - 6'b011011;
  /* TG68K_ALU.vhd:858:48  */
  assign n10966 = $unsigned(bs_shift) > $unsigned(6'b010001);
  /* TG68K_ALU.vhd:859:66  */
  assign n10968 = bs_shift - 6'b010010;
  /* TG68K_ALU.vhd:860:48  */
  assign n10970 = $unsigned(bs_shift) > $unsigned(6'b001000);
  /* TG68K_ALU.vhd:861:66  */
  assign n10972 = bs_shift - 6'b001001;
  /* TG68K_ALU.vhd:860:33  */
  assign n10973 = n10970 ? n10972 : bs_shift;
  /* TG68K_ALU.vhd:858:33  */
  assign n10974 = n10966 ? n10968 : n10973;
  /* TG68K_ALU.vhd:856:33  */
  assign n10975 = n10962 ? n10964 : n10974;
  /* TG68K_ALU.vhd:854:33  */
  assign n10976 = n10958 ? n10960 : n10975;
  /* TG68K_ALU.vhd:852:33  */
  assign n10977 = n10954 ? n10956 : n10976;
  /* TG68K_ALU.vhd:850:33  */
  assign n10978 = n10950 ? n10952 : n10977;
  /* TG68K_ALU.vhd:848:33  */
  assign n10980 = n10948 ? 6'b000000 : n10978;
  /* TG68K_ALU.vhd:847:25  */
  assign n10982 = ring == 6'b001001;
  /* TG68K_ALU.vhd:866:45  */
  assign n10984 = $unsigned(bs_shift) > $unsigned(6'b110010);
  /* TG68K_ALU.vhd:867:66  */
  assign n10986 = bs_shift - 6'b110011;
  /* TG68K_ALU.vhd:868:48  */
  assign n10988 = $unsigned(bs_shift) > $unsigned(6'b100001);
  /* TG68K_ALU.vhd:869:66  */
  assign n10990 = bs_shift - 6'b100010;
  /* TG68K_ALU.vhd:870:48  */
  assign n10992 = $unsigned(bs_shift) > $unsigned(6'b010000);
  /* TG68K_ALU.vhd:871:66  */
  assign n10994 = bs_shift - 6'b010001;
  /* TG68K_ALU.vhd:870:33  */
  assign n10995 = n10992 ? n10994 : bs_shift;
  /* TG68K_ALU.vhd:868:33  */
  assign n10996 = n10988 ? n10990 : n10995;
  /* TG68K_ALU.vhd:866:33  */
  assign n10997 = n10984 ? n10986 : n10996;
  /* TG68K_ALU.vhd:865:25  */
  assign n10999 = ring == 6'b010001;
  /* TG68K_ALU.vhd:876:45  */
  assign n11001 = $unsigned(bs_shift) > $unsigned(6'b100000);
  /* TG68K_ALU.vhd:877:66  */
  assign n11003 = bs_shift - 6'b100001;
  /* TG68K_ALU.vhd:876:33  */
  assign n11004 = n11001 ? n11003 : bs_shift;
  /* TG68K_ALU.vhd:875:25  */
  assign n11006 = ring == 6'b100001;
  /* TG68K_ALU.vhd:881:74  */
  assign n11007 = bs_shift[2:0]; // extract
  /* TG68K_ALU.vhd:881:64  */
  assign n11009 = {3'b000, n11007};
  /* TG68K_ALU.vhd:881:25  */
  assign n11011 = ring == 6'b001000;
  /* TG68K_ALU.vhd:882:74  */
  assign n11012 = bs_shift[3:0]; // extract
  /* TG68K_ALU.vhd:882:64  */
  assign n11014 = {2'b00, n11012};
  /* TG68K_ALU.vhd:882:25  */
  assign n11016 = ring == 6'b010000;
  /* TG68K_ALU.vhd:883:74  */
  assign n11017 = bs_shift[4:0]; // extract
  /* TG68K_ALU.vhd:883:64  */
  assign n11019 = {1'b0, n11017};
  /* TG68K_ALU.vhd:883:25  */
  assign n11021 = ring == 6'b100000;
  assign n11022 = {n11021, n11016, n11011, n11006, n10999, n10982};
  /* TG68K_ALU.vhd:846:17  */
  always @*
    case (n11022)
      6'b100000: n11024 = n11019;
      6'b010000: n11024 = n11014;
      6'b001000: n11024 = n11009;
      6'b000100: n11024 = n11004;
      6'b000010: n11024 = n10997;
      6'b000001: n11024 = n10980;
      default: n11024 = 6'b000000;
    endcase
  /* TG68K_ALU.vhd:888:30  */
  assign n11025 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:888:33  */
  assign n11026 = ~n11025;
  /* TG68K_ALU.vhd:889:39  */
  assign n11027 = ring - bs_shift_mod;
  /* TG68K_ALU.vhd:888:17  */
  assign n11028 = n11026 ? n11027 : bs_shift_mod;
  /* TG68K_ALU.vhd:891:28  */
  assign n11029 = rot_bits[1]; // extract
  /* TG68K_ALU.vhd:891:31  */
  assign n11030 = ~n11029;
  /* TG68K_ALU.vhd:892:38  */
  assign n11031 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:892:41  */
  assign n11032 = ~n11031;
  /* TG68K_ALU.vhd:893:45  */
  assign n11034 = 6'b100000 - bs_shift_mod;
  /* TG68K_ALU.vhd:892:25  */
  assign n11035 = n11032 ? n11034 : n11028;
  /* TG68K_ALU.vhd:895:37  */
  assign n11036 = bs_shift == ring;
  /* TG68K_ALU.vhd:896:46  */
  assign n11037 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:896:49  */
  assign n11038 = ~n11037;
  /* TG68K_ALU.vhd:897:53  */
  assign n11040 = 6'b100000 - ring;
  /* TG68K_ALU.vhd:896:33  */
  assign n11041 = n11038 ? n11040 : ring;
  /* TG68K_ALU.vhd:895:25  */
  assign n11042 = n11036 ? n11041 : n11035;
  /* TG68K_ALU.vhd:902:37  */
  assign n11043 = $unsigned(bs_shift) > $unsigned(ring);
  /* TG68K_ALU.vhd:903:46  */
  assign n11044 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:903:49  */
  assign n11045 = ~n11044;
  /* TG68K_ALU.vhd:907:55  */
  assign n11047 = ring + 6'b000001;
  /* TG68K_ALU.vhd:903:33  */
  assign n11049 = n11045 ? 6'b000000 : n11047;
  /* TG68K_ALU.vhd:891:17  */
  assign n11051 = n11055 ? 1'b0 : n10945;
  /* TG68K_ALU.vhd:902:25  */
  assign n11052 = n11043 ? n11049 : n11042;
  /* TG68K_ALU.vhd:902:25  */
  assign n11053 = n11045 & n11043;
  /* TG68K_ALU.vhd:891:17  */
  assign n11054 = n11030 ? n11052 : n11028;
  /* TG68K_ALU.vhd:891:17  */
  assign n11055 = n11053 & n11030;
  /* TG68K_ALU.vhd:915:50  */
  assign n11056 = asr_sign[31:0]; // extract
  /* TG68K_ALU.vhd:915:74  */
  assign n11057 = hot_msb[31:0]; // extract
  /* TG68K_ALU.vhd:915:64  */
  assign n11058 = n11056 | n11057;
  assign n11060 = n11059[0]; // extract
  /* TG68K_ALU.vhd:916:28  */
  assign n11062 = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:916:48  */
  assign n11063 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:916:51  */
  assign n11064 = ~n11063;
  /* TG68K_ALU.vhd:916:34  */
  assign n11065 = n11064 & n11062;
  /* TG68K_ALU.vhd:916:56  */
  assign n11066 = msb & n11065;
  /* TG68K_ALU.vhd:917:49  */
  assign n11067 = asr_sign[32:1]; // extract
  /* TG68K_ALU.vhd:917:38  */
  assign n11068 = alu | n11067;
  /* TG68K_ALU.vhd:918:37  */
  assign n11069 = $unsigned(bs_shift) > $unsigned(ring);
  /* TG68K_ALU.vhd:916:17  */
  assign n11071 = n11073 ? 1'b1 : n11051;
  /* TG68K_ALU.vhd:916:17  */
  assign n11072 = n11066 ? n11068 : alu;
  /* TG68K_ALU.vhd:916:17  */
  assign n11073 = n11069 & n11066;
  /* TG68K_ALU.vhd:923:43  */
  assign n11075 = {1'b0, op1out};
  /* TG68K_ALU.vhd:924:32  */
  assign n11076 = exe_opcode[7:6]; // extract
  /* TG68K_ALU.vhd:926:46  */
  assign n11077 = op1out[7]; // extract
  /* TG68K_ALU.vhd:929:44  */
  assign n11081 = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:930:59  */
  assign n11082 = n11806[4]; // extract
  assign n11083 = n11078[0]; // extract
  /* TG68K_ALU.vhd:929:33  */
  assign n11084 = n11081 ? n11082 : n11083;
  assign n11085 = n11078[23:1]; // extract
  /* TG68K_ALU.vhd:925:25  */
  assign n11087 = n11076 == 2'b00;
  /* TG68K_ALU.vhd:933:46  */
  assign n11088 = op1out[15]; // extract
  /* TG68K_ALU.vhd:936:44  */
  assign n11092 = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:937:60  */
  assign n11093 = n11806[4]; // extract
  assign n11094 = n11089[0]; // extract
  /* TG68K_ALU.vhd:936:33  */
  assign n11095 = n11092 ? n11093 : n11094;
  assign n11096 = n11089[15:1]; // extract
  /* TG68K_ALU.vhd:932:25  */
  assign n11098 = n11076 == 2'b01;
  /* TG68K_ALU.vhd:932:34  */
  assign n11100 = n11076 == 2'b11;
  /* TG68K_ALU.vhd:932:34  */
  assign n11101 = n11098 | n11100;
  /* TG68K_ALU.vhd:940:46  */
  assign n11102 = op1out[31]; // extract
  /* TG68K_ALU.vhd:941:44  */
  assign n11104 = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:942:60  */
  assign n11105 = n11806[4]; // extract
  assign n11106 = n11075[32]; // extract
  /* TG68K_ALU.vhd:941:33  */
  assign n11107 = n11104 ? n11105 : n11106;
  /* TG68K_ALU.vhd:939:25  */
  assign n11109 = n11076 == 2'b10;
  assign n11110 = {n11109, n11101, n11087};
  assign n11111 = n11075[8]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11112 = n11111;
      3'b010: n11112 = n11111;
      3'b001: n11112 = n11084;
      default: n11112 = n11111;
    endcase
  assign n11113 = n11085[6:0]; // extract
  assign n11114 = n11075[15:9]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11115 = n11114;
      3'b010: n11115 = n11114;
      3'b001: n11115 = n11113;
      default: n11115 = n11114;
    endcase
  assign n11116 = n11085[7]; // extract
  assign n11117 = n11075[16]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11118 = n11117;
      3'b010: n11118 = n11095;
      3'b001: n11118 = n11116;
      default: n11118 = n11117;
    endcase
  assign n11119 = n11085[22:8]; // extract
  assign n11120 = n11075[31:17]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11121 = n11120;
      3'b010: n11121 = n11096;
      3'b001: n11121 = n11119;
      default: n11121 = n11120;
    endcase
  assign n11122 = n11075[32]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11123 = n11107;
      3'b010: n11123 = n11122;
      3'b001: n11123 = n11122;
      default: n11123 = n11122;
    endcase
  assign n11125 = n11075[7:0]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11129 = n11102;
      3'b010: n11129 = n11088;
      3'b001: n11129 = n11077;
      default: n11129 = msb;
    endcase
  assign n11130 = n11079[7:0]; // extract
  assign n11131 = n11072[15:8]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11132 = n11131;
      3'b010: n11132 = n11131;
      3'b001: n11132 = n11130;
      default: n11132 = n11131;
    endcase
  assign n11133 = n11079[23:8]; // extract
  assign n11134 = n11072[31:16]; // extract
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n11110)
      3'b100: n11135 = n11134;
      3'b010: n11135 = 16'b0000000000000000;
      3'b001: n11135 = n11133;
      default: n11135 = n11134;
    endcase
  assign n11137 = n11072[7:0]; // extract
  /* TG68K_ALU.vhd:946:71  */
  assign n11139 = {33'b000000000000000000000000000000000, vector};
  /* TG68K_ALU.vhd:946:84  */
  assign n11140 = {25'b0, bit_nr};  //  uext
  /* TG68K_ALU.vhd:946:80  */
  assign n11141 = {1'b0, n11140};  //  uext
  /* TG68K_ALU.vhd:946:80  */
  assign n11142 = n11139 << n11141;
  /* TG68K_ALU.vhd:957:24  */
  assign n11146 = exec[17]; // extract
  /* TG68K_ALU.vhd:958:58  */
  assign n11147 = last_data_read[7:0]; // extract
  /* TG68K_ALU.vhd:958:40  */
  assign n11148 = n11806 & n11147;
  /* TG68K_ALU.vhd:959:27  */
  assign n11149 = exec[18]; // extract
  /* TG68K_ALU.vhd:960:58  */
  assign n11150 = last_data_read[7:0]; // extract
  /* TG68K_ALU.vhd:960:40  */
  assign n11151 = n11806 ^ n11150;
  /* TG68K_ALU.vhd:961:27  */
  assign n11152 = exec[19]; // extract
  /* TG68K_ALU.vhd:962:57  */
  assign n11153 = last_data_read[7:0]; // extract
  /* TG68K_ALU.vhd:962:40  */
  assign n11154 = n11806 | n11153;
  /* TG68K_ALU.vhd:964:40  */
  assign n11155 = op2out[7:0]; // extract
  /* TG68K_ALU.vhd:961:17  */
  assign n11156 = n11152 ? n11154 : n11155;
  /* TG68K_ALU.vhd:959:17  */
  assign n11157 = n11149 ? n11151 : n11156;
  /* TG68K_ALU.vhd:957:17  */
  assign n11158 = n11146 ? n11148 : n11157;
  /* TG68K_ALU.vhd:971:24  */
  assign n11159 = exec[28]; // extract
  /* TG68K_ALU.vhd:971:50  */
  assign n11160 = n11806[2]; // extract
  /* TG68K_ALU.vhd:971:53  */
  assign n11161 = ~n11160;
  /* TG68K_ALU.vhd:971:41  */
  assign n11162 = n11161 & n11159;
  /* TG68K_ALU.vhd:973:28  */
  assign n11163 = op1in[7:0]; // extract
  /* TG68K_ALU.vhd:973:40  */
  assign n11165 = n11163 == 8'b00000000;
  /* TG68K_ALU.vhd:975:33  */
  assign n11167 = op1in[15:8]; // extract
  /* TG68K_ALU.vhd:975:46  */
  assign n11169 = n11167 == 8'b00000000;
  /* TG68K_ALU.vhd:977:41  */
  assign n11171 = op1in[31:16]; // extract
  /* TG68K_ALU.vhd:977:55  */
  assign n11173 = n11171 == 16'b0000000000000000;
  /* TG68K_ALU.vhd:977:33  */
  assign n11176 = n11173 ? 1'b1 : 1'b0;
  assign n11177 = {n11176, 1'b1};
  /* TG68K_ALU.vhd:975:25  */
  assign n11179 = n11169 ? n11177 : 2'b00;
  assign n11180 = {n11179, 1'b1};
  /* TG68K_ALU.vhd:973:17  */
  assign n11182 = n11165 ? n11180 : 3'b000;
  /* TG68K_ALU.vhd:971:17  */
  assign n11184 = n11162 ? 3'b000 : n11182;
  /* TG68K_ALU.vhd:984:32  */
  assign n11187 = exe_datatype == 2'b00;
  /* TG68K_ALU.vhd:985:43  */
  assign n11188 = op1in[7]; // extract
  /* TG68K_ALU.vhd:985:53  */
  assign n11189 = flag_z[0]; // extract
  /* TG68K_ALU.vhd:985:46  */
  assign n11190 = {n11188, n11189};
  /* TG68K_ALU.vhd:985:67  */
  assign n11191 = addsub_ofl[0]; // extract
  /* TG68K_ALU.vhd:985:56  */
  assign n11192 = {n11190, n11191};
  /* TG68K_ALU.vhd:985:76  */
  assign n11193 = n9689[0]; // extract
  /* TG68K_ALU.vhd:985:70  */
  assign n11194 = {n11192, n11193};
  /* TG68K_ALU.vhd:986:32  */
  assign n11195 = exec[12]; // extract
  /* TG68K_ALU.vhd:986:53  */
  assign n11196 = exec[13]; // extract
  /* TG68K_ALU.vhd:986:46  */
  assign n11197 = n11195 | n11196;
  assign n11198 = {vflag_a, bcd_a_carry};
  assign n11199 = n11194[1:0]; // extract
  /* TG68K_ALU.vhd:986:25  */
  assign n11200 = n11197 ? n11198 : n11199;
  assign n11201 = n11194[3:2]; // extract
  /* TG68K_ALU.vhd:990:35  */
  assign n11203 = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:990:48  */
  assign n11204 = exec[10]; // extract
  /* TG68K_ALU.vhd:990:41  */
  assign n11205 = n11203 | n11204;
  /* TG68K_ALU.vhd:991:43  */
  assign n11206 = op1in[31]; // extract
  /* TG68K_ALU.vhd:991:54  */
  assign n11207 = flag_z[2]; // extract
  /* TG68K_ALU.vhd:991:47  */
  assign n11208 = {n11206, n11207};
  /* TG68K_ALU.vhd:991:68  */
  assign n11209 = addsub_ofl[2]; // extract
  /* TG68K_ALU.vhd:991:57  */
  assign n11210 = {n11208, n11209};
  /* TG68K_ALU.vhd:991:77  */
  assign n11211 = n9689[2]; // extract
  /* TG68K_ALU.vhd:991:71  */
  assign n11212 = {n11210, n11211};
  /* TG68K_ALU.vhd:993:43  */
  assign n11213 = op1in[15]; // extract
  /* TG68K_ALU.vhd:993:54  */
  assign n11214 = flag_z[1]; // extract
  /* TG68K_ALU.vhd:993:47  */
  assign n11215 = {n11213, n11214};
  /* TG68K_ALU.vhd:993:68  */
  assign n11216 = addsub_ofl[1]; // extract
  /* TG68K_ALU.vhd:993:57  */
  assign n11217 = {n11215, n11216};
  /* TG68K_ALU.vhd:993:77  */
  assign n11218 = n9689[1]; // extract
  /* TG68K_ALU.vhd:993:71  */
  assign n11219 = {n11217, n11218};
  /* TG68K_ALU.vhd:990:17  */
  assign n11220 = n11205 ? n11212 : n11219;
  assign n11221 = {n11201, n11200};
  /* TG68K_ALU.vhd:984:17  */
  assign n11222 = n11187 ? n11221 : n11220;
  /* TG68K_ALU.vhd:1000:40  */
  assign n11224 = exec[59]; // extract
  /* TG68K_ALU.vhd:1000:55  */
  assign n11225 = n11224 | set_stop;
  /* TG68K_ALU.vhd:1001:71  */
  assign n11226 = data_read[7:0]; // extract
  /* TG68K_ALU.vhd:1000:33  */
  assign n11227 = n11225 ? n11226 : n11806;
  /* TG68K_ALU.vhd:1003:40  */
  assign n11228 = exec[60]; // extract
  /* TG68K_ALU.vhd:1004:71  */
  assign n11229 = data_read[7:0]; // extract
  /* TG68K_ALU.vhd:1003:33  */
  assign n11230 = n11228 ? n11229 : n11227;
  /* TG68K_ALU.vhd:1007:40  */
  assign n11231 = exec[9]; // extract
  /* TG68K_ALU.vhd:1007:66  */
  assign n11232 = ~decodeopc;
  /* TG68K_ALU.vhd:1007:53  */
  assign n11233 = n11232 & n11231;
  /* TG68K_ALU.vhd:1008:65  */
  assign n11234 = set_flags[3]; // extract
  /* TG68K_ALU.vhd:1008:69  */
  assign n11235 = n11234 ^ rot_rot;
  /* TG68K_ALU.vhd:1008:82  */
  assign n11236 = n11235 | asl_vflag;
  /* TG68K_ALU.vhd:1007:33  */
  assign n11238 = n11233 ? n11236 : 1'b0;
  /* TG68K_ALU.vhd:1012:40  */
  assign n11239 = exec[51]; // extract
  /* TG68K_ALU.vhd:1015:56  */
  assign n11241 = micro_state == 7'b0110011;
  /* TG68K_ALU.vhd:1017:62  */
  assign n11242 = exe_opcode[8]; // extract
  /* TG68K_ALU.vhd:1017:65  */
  assign n11243 = ~n11242;
  /* TG68K_ALU.vhd:1019:92  */
  assign n11244 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1019:82  */
  assign n11245 = ~n11244;
  /* TG68K_ALU.vhd:1019:81  */
  assign n11247 = {1'b0, n11245};
  /* TG68K_ALU.vhd:1019:96  */
  assign n11249 = {n11247, 2'b00};
  /* TG68K_ALU.vhd:1017:49  */
  assign n11251 = n11243 ? n11249 : 4'b0100;
  assign n11252 = n11230[3:0]; // extract
  /* TG68K_ALU.vhd:1015:41  */
  assign n11253 = n11241 ? n11251 : n11252;
  /* TG68K_ALU.vhd:1024:43  */
  assign n11254 = exec[49]; // extract
  /* TG68K_ALU.vhd:1024:53  */
  assign n11255 = ~n11254;
  /* TG68K_ALU.vhd:1025:61  */
  assign n11256 = n11806[3:0]; // extract
  /* TG68K_ALU.vhd:1026:48  */
  assign n11257 = exec[3]; // extract
  /* TG68K_ALU.vhd:1027:70  */
  assign n11258 = set_flags[0]; // extract
  /* TG68K_ALU.vhd:1028:51  */
  assign n11259 = exec[9]; // extract
  /* TG68K_ALU.vhd:1028:76  */
  assign n11261 = rot_bits != 2'b11;
  /* TG68K_ALU.vhd:1028:64  */
  assign n11262 = n11261 & n11259;
  /* TG68K_ALU.vhd:1028:91  */
  assign n11263 = exec[23]; // extract
  /* TG68K_ALU.vhd:1028:100  */
  assign n11264 = ~n11263;
  /* TG68K_ALU.vhd:1028:83  */
  assign n11265 = n11264 & n11262;
  /* TG68K_ALU.vhd:1030:51  */
  assign n11266 = exec[81]; // extract
  assign n11267 = n11230[4]; // extract
  /* TG68K_ALU.vhd:1030:41  */
  assign n11268 = n11266 ? bs_x : n11267;
  /* TG68K_ALU.vhd:1028:41  */
  assign n11269 = n11265 ? rot_x : n11268;
  /* TG68K_ALU.vhd:1026:41  */
  assign n11270 = n11257 ? n11258 : n11269;
  /* TG68K_ALU.vhd:1034:49  */
  assign n11271 = exec[8]; // extract
  /* TG68K_ALU.vhd:1034:65  */
  assign n11272 = exec[86]; // extract
  /* TG68K_ALU.vhd:1034:58  */
  assign n11273 = n11271 | n11272;
  /* TG68K_ALU.vhd:1036:51  */
  assign n11274 = exec[21]; // extract
  /* TG68K_ALU.vhd:1036:65  */
  assign n11276 = 1'b1 & n11274;
  /* TG68K_ALU.vhd:1039:65  */
  assign n11278 = exe_opcode[15]; // extract
  /* TG68K_ALU.vhd:1039:74  */
  assign n11280 = n11278 | 1'b0;
  /* TG68K_ALU.vhd:1040:83  */
  assign n11281 = op1in[15]; // extract
  /* TG68K_ALU.vhd:1040:94  */
  assign n11282 = flag_z[1]; // extract
  /* TG68K_ALU.vhd:1040:87  */
  assign n11283 = {n11281, n11282};
  /* TG68K_ALU.vhd:1040:97  */
  assign n11285 = {n11283, 2'b00};
  /* TG68K_ALU.vhd:1042:83  */
  assign n11286 = op1in[31]; // extract
  /* TG68K_ALU.vhd:1042:94  */
  assign n11287 = flag_z[2]; // extract
  /* TG68K_ALU.vhd:1042:87  */
  assign n11288 = {n11286, n11287};
  /* TG68K_ALU.vhd:1042:97  */
  assign n11290 = {n11288, 2'b00};
  /* TG68K_ALU.vhd:1039:49  */
  assign n11291 = n11280 ? n11285 : n11290;
  /* TG68K_ALU.vhd:1037:49  */
  assign n11292 = v_flag ? 4'b1010 : n11291;
  /* TG68K_ALU.vhd:1044:51  */
  assign n11293 = exec[68]; // extract
  /* TG68K_ALU.vhd:1044:72  */
  assign n11295 = 1'b1 & n11293;
  /* TG68K_ALU.vhd:1045:70  */
  assign n11296 = set_flags[3]; // extract
  /* TG68K_ALU.vhd:1046:70  */
  assign n11297 = set_flags[2]; // extract
  /* TG68K_ALU.vhd:1046:83  */
  assign n11298 = n11806[2]; // extract
  /* TG68K_ALU.vhd:1046:74  */
  assign n11299 = n11297 & n11298;
  /* TG68K_ALU.vhd:1049:51  */
  assign n11302 = exec[67]; // extract
  /* TG68K_ALU.vhd:1049:71  */
  assign n11304 = 1'b1 & n11302;
  /* TG68K_ALU.vhd:1050:70  */
  assign n11305 = set_flags[3]; // extract
  /* TG68K_ALU.vhd:1051:70  */
  assign n11306 = set_flags[2]; // extract
  /* TG68K_ALU.vhd:1054:51  */
  assign n11308 = exec[5]; // extract
  /* TG68K_ALU.vhd:1054:70  */
  assign n11309 = exec[6]; // extract
  /* TG68K_ALU.vhd:1054:63  */
  assign n11310 = n11308 | n11309;
  /* TG68K_ALU.vhd:1054:90  */
  assign n11311 = exec[7]; // extract
  /* TG68K_ALU.vhd:1054:83  */
  assign n11312 = n11310 | n11311;
  /* TG68K_ALU.vhd:1054:110  */
  assign n11313 = exec[0]; // extract
  /* TG68K_ALU.vhd:1054:103  */
  assign n11314 = n11312 | n11313;
  /* TG68K_ALU.vhd:1054:131  */
  assign n11315 = exec[1]; // extract
  /* TG68K_ALU.vhd:1054:124  */
  assign n11316 = n11314 | n11315;
  /* TG68K_ALU.vhd:1054:153  */
  assign n11317 = exec[15]; // extract
  /* TG68K_ALU.vhd:1054:146  */
  assign n11318 = n11316 | n11317;
  /* TG68K_ALU.vhd:1054:174  */
  assign n11319 = exec[75]; // extract
  /* TG68K_ALU.vhd:1054:167  */
  assign n11320 = n11318 | n11319;
  /* TG68K_ALU.vhd:1054:194  */
  assign n11321 = exec[20]; // extract
  /* TG68K_ALU.vhd:1054:208  */
  assign n11323 = 1'b1 & n11321;
  /* TG68K_ALU.vhd:1054:186  */
  assign n11324 = n11320 | n11323;
  /* TG68K_ALU.vhd:1057:56  */
  assign n11327 = exec[75]; // extract
  assign n11328 = set_flags[3]; // extract
  /* TG68K_ALU.vhd:1057:49  */
  assign n11329 = n11327 ? bf_nflag : n11328;
  assign n11330 = set_flags[2]; // extract
  /* TG68K_ALU.vhd:1060:51  */
  assign n11331 = exec[9]; // extract
  /* TG68K_ALU.vhd:1061:79  */
  assign n11332 = set_flags[3:2]; // extract
  /* TG68K_ALU.vhd:1063:60  */
  assign n11334 = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:1063:81  */
  assign n11335 = set_flags[3]; // extract
  /* TG68K_ALU.vhd:1063:85  */
  assign n11336 = n11335 ^ rot_rot;
  /* TG68K_ALU.vhd:1063:98  */
  assign n11337 = n11336 | asl_vflag;
  /* TG68K_ALU.vhd:1063:66  */
  assign n11338 = n11337 & n11334;
  /* TG68K_ALU.vhd:1063:49  */
  assign n11341 = n11338 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1068:51  */
  assign n11342 = exec[81]; // extract
  /* TG68K_ALU.vhd:1069:79  */
  assign n11343 = set_flags[3:2]; // extract
  /* TG68K_ALU.vhd:1072:51  */
  assign n11344 = exec[14]; // extract
  /* TG68K_ALU.vhd:1073:61  */
  assign n11345 = ~one_bit_in;
  /* TG68K_ALU.vhd:1074:51  */
  assign n11346 = exec[87]; // extract
  /* TG68K_ALU.vhd:1079:63  */
  assign n11347 = last_flags1[0]; // extract
  /* TG68K_ALU.vhd:1079:66  */
  assign n11348 = ~n11347;
  /* TG68K_ALU.vhd:1080:74  */
  assign n11349 = n11806[0]; // extract
  /* TG68K_ALU.vhd:1080:95  */
  assign n11350 = set_flags[0]; // extract
  /* TG68K_ALU.vhd:1080:82  */
  assign n11351 = ~n11350;
  /* TG68K_ALU.vhd:1080:116  */
  assign n11352 = set_flags[2]; // extract
  /* TG68K_ALU.vhd:1080:103  */
  assign n11353 = ~n11352;
  /* TG68K_ALU.vhd:1080:99  */
  assign n11354 = n11351 & n11353;
  /* TG68K_ALU.vhd:1080:78  */
  assign n11355 = n11349 | n11354;
  /* TG68K_ALU.vhd:1082:75  */
  assign n11356 = n11806[0]; // extract
  /* TG68K_ALU.vhd:1082:92  */
  assign n11357 = set_flags[0]; // extract
  /* TG68K_ALU.vhd:1082:79  */
  assign n11358 = n11356 ^ n11357;
  /* TG68K_ALU.vhd:1082:111  */
  assign n11359 = n11806[2]; // extract
  /* TG68K_ALU.vhd:1082:102  */
  assign n11360 = ~n11359;
  /* TG68K_ALU.vhd:1082:97  */
  assign n11361 = n11358 & n11360;
  /* TG68K_ALU.vhd:1082:132  */
  assign n11362 = set_flags[2]; // extract
  /* TG68K_ALU.vhd:1082:119  */
  assign n11363 = ~n11362;
  /* TG68K_ALU.vhd:1082:115  */
  assign n11364 = n11361 & n11363;
  /* TG68K_ALU.vhd:1079:49  */
  assign n11365 = n11348 ? n11355 : n11364;
  /* TG68K_ALU.vhd:1085:66  */
  assign n11367 = n11806[2]; // extract
  /* TG68K_ALU.vhd:1085:82  */
  assign n11368 = set_flags[2]; // extract
  /* TG68K_ALU.vhd:1085:70  */
  assign n11369 = n11367 | n11368;
  /* TG68K_ALU.vhd:1086:76  */
  assign n11370 = last_flags1[0]; // extract
  /* TG68K_ALU.vhd:1086:61  */
  assign n11371 = ~n11370;
  /* TG68K_ALU.vhd:1087:51  */
  assign n11372 = exec[31]; // extract
  /* TG68K_ALU.vhd:1088:64  */
  assign n11374 = exe_datatype == 2'b01;
  /* TG68K_ALU.vhd:1089:75  */
  assign n11375 = op1out[15]; // extract
  /* TG68K_ALU.vhd:1091:75  */
  assign n11376 = op1out[31]; // extract
  /* TG68K_ALU.vhd:1088:49  */
  assign n11377 = n11374 ? n11375 : n11376;
  /* TG68K_ALU.vhd:1093:58  */
  assign n11378 = op1out[15:0]; // extract
  /* TG68K_ALU.vhd:1093:71  */
  assign n11380 = n11378 == 16'b0000000000000000;
  /* TG68K_ALU.vhd:1093:97  */
  assign n11382 = exe_datatype == 2'b01;
  /* TG68K_ALU.vhd:1093:112  */
  assign n11383 = op1out[31:16]; // extract
  /* TG68K_ALU.vhd:1093:126  */
  assign n11385 = n11383 == 16'b0000000000000000;
  /* TG68K_ALU.vhd:1093:103  */
  assign n11386 = n11382 | n11385;
  /* TG68K_ALU.vhd:1093:80  */
  assign n11387 = n11386 & n11380;
  /* TG68K_ALU.vhd:1093:49  */
  assign n11390 = n11387 ? 1'b1 : 1'b0;
  assign n11393 = {n11377, n11390, 1'b0, 1'b0};
  assign n11394 = n11230[3:0]; // extract
  /* TG68K_ALU.vhd:1087:41  */
  assign n11395 = n11372 ? n11393 : n11394;
  assign n11396 = {n11371, n11369, 1'b0, n11365};
  /* TG68K_ALU.vhd:1074:41  */
  assign n11397 = n11346 ? n11396 : n11395;
  assign n11398 = n11397[1:0]; // extract
  assign n11399 = n11230[1:0]; // extract
  /* TG68K_ALU.vhd:1072:41  */
  assign n11400 = n11344 ? n11399 : n11398;
  assign n11401 = n11397[2]; // extract
  /* TG68K_ALU.vhd:1072:41  */
  assign n11402 = n11344 ? n11345 : n11401;
  assign n11403 = n11397[3]; // extract
  assign n11404 = n11230[3]; // extract
  /* TG68K_ALU.vhd:1072:41  */
  assign n11405 = n11344 ? n11404 : n11403;
  assign n11406 = {n11405, n11402, n11400};
  assign n11407 = {n11343, bs_v, bs_c};
  /* TG68K_ALU.vhd:1068:41  */
  assign n11408 = n11342 ? n11407 : n11406;
  assign n11409 = {n11332, n11341, rot_c};
  /* TG68K_ALU.vhd:1060:41  */
  assign n11410 = n11331 ? n11409 : n11408;
  assign n11411 = {n11329, n11330, 2'b00};
  /* TG68K_ALU.vhd:1054:41  */
  assign n11412 = n11324 ? n11411 : n11410;
  assign n11413 = {n11305, n11306, set_mv_flag, 1'b0};
  /* TG68K_ALU.vhd:1049:41  */
  assign n11414 = n11304 ? n11413 : n11412;
  assign n11415 = {n11296, n11299, 1'b0, 1'b0};
  /* TG68K_ALU.vhd:1044:41  */
  assign n11416 = n11295 ? n11415 : n11414;
  /* TG68K_ALU.vhd:1036:41  */
  assign n11417 = n11276 ? n11292 : n11416;
  /* TG68K_ALU.vhd:1034:41  */
  assign n11418 = n11273 ? set_flags : n11417;
  assign n11419 = {n11270, n11418};
  assign n11420 = n11230[4:0]; // extract
  /* TG68K_ALU.vhd:1024:33  */
  assign n11421 = n11255 ? n11419 : n11420;
  /* TG68K_ALU.vhd:1024:33  */
  assign n11422 = n11255 ? n11256 : last_flags1;
  assign n11423 = n11421[3:0]; // extract
  /* TG68K_ALU.vhd:1014:33  */
  assign n11424 = z_error ? n11253 : n11423;
  assign n11425 = n11421[4]; // extract
  assign n11426 = n11230[4]; // extract
  /* TG68K_ALU.vhd:1014:33  */
  assign n11427 = z_error ? n11426 : n11425;
  /* TG68K_ALU.vhd:1014:33  */
  assign n11428 = z_error ? last_flags1 : n11422;
  assign n11429 = {n11427, n11424};
  assign n11430 = ccrin[4:0]; // extract
  /* TG68K_ALU.vhd:1012:33  */
  assign n11431 = n11239 ? n11430 : n11429;
  assign n11432 = ccrin[7:5]; // extract
  assign n11433 = n11230[7:5]; // extract
  /* TG68K_ALU.vhd:1012:33  */
  assign n11434 = n11239 ? n11432 : n11433;
  /* TG68K_ALU.vhd:1012:33  */
  assign n11436 = n11239 ? last_flags1 : n11428;
  assign n11437 = {n11434, n11431};
  /* TG68K_ALU.vhd:999:25  */
  assign n11438 = clkena_lw ? n11437 : n11806;
  /* TG68K_ALU.vhd:999:25  */
  assign n11439 = clkena_lw ? n11436 : last_flags1;
  /* TG68K_ALU.vhd:999:25  */
  assign n11440 = clkena_lw ? n11238 : asl_vflag;
  /* TG68K_ALU.vhd:997:25  */
  assign n11442 = reset ? 8'b00000000 : n11438;
  /* TG68K_ALU.vhd:997:25  */
  assign n11443 = reset ? last_flags1 : n11439;
  /* TG68K_ALU.vhd:997:25  */
  assign n11444 = reset ? asl_vflag : n11440;
  assign n11446 = n11442[4:0]; // extract
  assign n11447 = {3'b000, n11446};
  /* TG68K_ALU.vhd:1128:38  */
  assign n11454 = exe_opcode[15]; // extract
  /* TG68K_ALU.vhd:1129:59  */
  assign n11455 = reg_qa[15]; // extract
  /* TG68K_ALU.vhd:1129:49  */
  assign n11456 = n11455 & signedop;
  /* TG68K_ALU.vhd:1129:33  */
  assign n11459 = n11456 ? 32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
  /* TG68K_ALU.vhd:1134:59  */
  assign n11460 = op2out[15]; // extract
  /* TG68K_ALU.vhd:1134:49  */
  assign n11461 = n11460 & signedop;
  /* TG68K_ALU.vhd:1134:33  */
  assign n11464 = n11461 ? 32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
  /* TG68K_ALU.vhd:1140:63  */
  assign n11465 = reg_qa[31:16]; // extract
  /* TG68K_ALU.vhd:1141:63  */
  assign n11466 = op2out[31:16]; // extract
  /* TG68K_ALU.vhd:1142:59  */
  assign n11467 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1142:49  */
  assign n11468 = n11467 & signedop;
  /* TG68K_ALU.vhd:1142:33  */
  assign n11471 = n11468 ? 16'b1111111111111111 : 16'b0000000000000000;
  /* TG68K_ALU.vhd:1147:59  */
  assign n11472 = op2out[31]; // extract
  /* TG68K_ALU.vhd:1147:49  */
  assign n11473 = n11472 & signedop;
  /* TG68K_ALU.vhd:1147:33  */
  assign n11476 = n11473 ? 16'b1111111111111111 : 16'b0000000000000000;
  assign n11477 = {n11471, n11465};
  /* TG68K_ALU.vhd:1128:25  */
  assign n11478 = n11454 ? n11459 : n11477;
  assign n11479 = {n11476, n11466};
  /* TG68K_ALU.vhd:1128:25  */
  assign n11480 = n11454 ? n11464 : n11479;
  /* TG68K_ALU.vhd:1153:62  */
  assign n11481 = faktora[31:16]; // extract
  /* TG68K_ALU.vhd:1153:77  */
  assign n11482 = {n11481, faktora};
  /* TG68K_ALU.vhd:1153:108  */
  assign n11483 = reg_qa[15:0]; // extract
  /* TG68K_ALU.vhd:1153:100  */
  assign n11484 = {n11482, n11483};
  /* TG68K_ALU.vhd:1153:133  */
  assign n11485 = faktorb[31:16]; // extract
  /* TG68K_ALU.vhd:1153:148  */
  assign n11486 = {n11485, faktorb};
  /* TG68K_ALU.vhd:1153:179  */
  assign n11487 = op2out[15:0]; // extract
  /* TG68K_ALU.vhd:1153:171  */
  assign n11488 = {n11486, n11487};
  /* TG68K_ALU.vhd:1153:123  */
  assign n11489 = {64'b0, n11484};  //  uext
  /* TG68K_ALU.vhd:1153:123  */
  assign n11490 = {64'b0, n11488};  //  uext
  /* TG68K_ALU.vhd:1153:123  */
  assign n11491 = n11489 * n11490; // umul
  /* TG68K_ALU.vhd:1201:32  */
  assign n11492 = result_mulu[63:32]; // extract
  /* TG68K_ALU.vhd:1201:46  */
  assign n11494 = n11492 == 32'b00000000000000000000000000000000;
  /* TG68K_ALU.vhd:1201:72  */
  assign n11495 = ~signedop;
  /* TG68K_ALU.vhd:1201:91  */
  assign n11496 = result_mulu[31]; // extract
  /* TG68K_ALU.vhd:1201:95  */
  assign n11497 = ~n11496;
  /* TG68K_ALU.vhd:1201:77  */
  assign n11498 = n11495 | n11497;
  /* TG68K_ALU.vhd:1201:59  */
  assign n11499 = n11498 & n11494;
  /* TG68K_ALU.vhd:1202:37  */
  assign n11500 = result_mulu[63:32]; // extract
  /* TG68K_ALU.vhd:1202:51  */
  assign n11502 = n11500 == 32'b11111111111111111111111111111111;
  /* TG68K_ALU.vhd:1202:64  */
  assign n11503 = signedop & n11502;
  /* TG68K_ALU.vhd:1202:96  */
  assign n11504 = result_mulu[31]; // extract
  /* TG68K_ALU.vhd:1202:81  */
  assign n11505 = n11504 & n11503;
  /* TG68K_ALU.vhd:1201:102  */
  assign n11506 = n11499 | n11505;
  /* TG68K_ALU.vhd:1201:17  */
  assign n11509 = n11506 ? 1'b0 : 1'b1;
  /* TG68K_ALU.vhd:1227:77  */
  assign n11514 = result_mulu[63:32]; // extract
  /* TG68K_ALU.vhd:1240:32  */
  assign n11522 = opcode[15]; // extract
  /* TG68K_ALU.vhd:1240:47  */
  assign n11523 = opcode[8]; // extract
  /* TG68K_ALU.vhd:1240:37  */
  assign n11524 = n11522 & n11523;
  /* TG68K_ALU.vhd:1240:66  */
  assign n11525 = opcode[15]; // extract
  /* TG68K_ALU.vhd:1240:56  */
  assign n11526 = ~n11525;
  /* TG68K_ALU.vhd:1240:81  */
  assign n11527 = sndopc[11]; // extract
  /* TG68K_ALU.vhd:1240:71  */
  assign n11528 = n11526 & n11527;
  /* TG68K_ALU.vhd:1240:52  */
  assign n11529 = n11524 | n11528;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11531 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11532 = divs & n11531;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11533 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11534 = divs & n11533;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11535 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11536 = divs & n11535;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11537 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11538 = divs & n11537;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11539 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11540 = divs & n11539;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11541 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11542 = divs & n11541;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11543 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11544 = divs & n11543;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11545 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11546 = divs & n11545;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11547 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11548 = divs & n11547;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11549 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11550 = divs & n11549;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11551 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11552 = divs & n11551;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11553 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11554 = divs & n11553;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11555 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11556 = divs & n11555;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11557 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11558 = divs & n11557;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11559 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11560 = divs & n11559;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11561 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11562 = divs & n11561;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11563 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11564 = divs & n11563;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11565 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11566 = divs & n11565;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11567 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11568 = divs & n11567;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11569 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11570 = divs & n11569;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11571 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11572 = divs & n11571;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11573 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11574 = divs & n11573;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11575 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11576 = divs & n11575;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11577 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11578 = divs & n11577;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11579 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11580 = divs & n11579;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11581 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11582 = divs & n11581;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11583 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11584 = divs & n11583;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11585 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11586 = divs & n11585;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11587 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11588 = divs & n11587;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11589 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11590 = divs & n11589;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11591 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11592 = divs & n11591;
  /* TG68K_ALU.vhd:1242:68  */
  assign n11593 = reg_qa[31]; // extract
  /* TG68K_ALU.vhd:1242:58  */
  assign n11594 = divs & n11593;
  assign n11595 = {n11532, n11534, n11536, n11538};
  assign n11596 = {n11540, n11542, n11544, n11546};
  assign n11597 = {n11548, n11550, n11552, n11554};
  assign n11598 = {n11556, n11558, n11560, n11562};
  assign n11599 = {n11564, n11566, n11568, n11570};
  assign n11600 = {n11572, n11574, n11576, n11578};
  assign n11601 = {n11580, n11582, n11584, n11586};
  assign n11602 = {n11588, n11590, n11592, n11594};
  assign n11603 = {n11595, n11596, n11597, n11598};
  assign n11604 = {n11599, n11600, n11601, n11602};
  assign n11605 = {n11603, n11604};
  /* TG68K_ALU.vhd:1243:30  */
  assign n11606 = exe_opcode[15]; // extract
  /* TG68K_ALU.vhd:1243:39  */
  assign n11608 = n11606 | 1'b0;
  /* TG68K_ALU.vhd:1245:52  */
  assign n11609 = result_div_pre[15]; // extract
  /* TG68K_ALU.vhd:1248:38  */
  assign n11610 = exe_opcode[14]; // extract
  /* TG68K_ALU.vhd:1248:57  */
  assign n11611 = sndopc[10]; // extract
  /* TG68K_ALU.vhd:1248:47  */
  assign n11612 = n11611 & n11610;
  /* TG68K_ALU.vhd:1248:25  */
  assign n11613 = n11612 ? reg_qb : n11605;
  /* TG68K_ALU.vhd:1251:52  */
  assign n11614 = result_div_pre[31]; // extract
  /* TG68K_ALU.vhd:1243:17  */
  assign n11615 = n11608 ? n11609 : n11614;
  assign n11616 = {n11613, reg_qa};
  assign n11617 = n11616[15:0]; // extract
  /* TG68K_ALU.vhd:1243:17  */
  assign n11618 = n11608 ? 16'b0000000000000000 : n11617;
  assign n11619 = n11616[47:16]; // extract
  /* TG68K_ALU.vhd:1243:17  */
  assign n11620 = n11608 ? reg_qa : n11619;
  assign n11621 = n11616[63:48]; // extract
  assign n11622 = n11605[31:16]; // extract
  /* TG68K_ALU.vhd:1243:17  */
  assign n11623 = n11608 ? n11622 : n11621;
  /* TG68K_ALU.vhd:1253:42  */
  assign n11625 = opcode[15]; // extract
  /* TG68K_ALU.vhd:1253:46  */
  assign n11626 = ~n11625;
  /* TG68K_ALU.vhd:1253:33  */
  assign n11627 = signedop | n11626;
  /* TG68K_ALU.vhd:1254:44  */
  assign n11628 = op2out[31:16]; // extract
  /* TG68K_ALU.vhd:1253:17  */
  assign n11630 = n11627 ? n11628 : 16'b0000000000000000;
  /* TG68K_ALU.vhd:1258:43  */
  assign n11631 = op2out[31]; // extract
  /* TG68K_ALU.vhd:1258:33  */
  assign n11632 = n11631 & signedop;
  /* TG68K_ALU.vhd:1259:44  */
  assign n11633 = div_reg[63:31]; // extract
  /* TG68K_ALU.vhd:1259:64  */
  assign n11635 = {1'b1, op2out};
  /* TG68K_ALU.vhd:1259:59  */
  assign n11636 = n11633 + n11635;
  /* TG68K_ALU.vhd:1261:44  */
  assign n11637 = div_reg[63:31]; // extract
  /* TG68K_ALU.vhd:1261:64  */
  assign n11639 = {1'b0, op2outext};
  /* TG68K_ALU.vhd:1261:94  */
  assign n11640 = op2out[15:0]; // extract
  /* TG68K_ALU.vhd:1261:87  */
  assign n11641 = {n11639, n11640};
  /* TG68K_ALU.vhd:1261:59  */
  assign n11642 = n11637 - n11641;
  /* TG68K_ALU.vhd:1258:17  */
  assign n11643 = n11632 ? n11636 : n11642;
  /* TG68K_ALU.vhd:1266:43  */
  assign n11644 = div_sub[32]; // extract
  /* TG68K_ALU.vhd:1269:58  */
  assign n11645 = div_reg[62:31]; // extract
  /* TG68K_ALU.vhd:1271:58  */
  assign n11646 = div_sub[31:0]; // extract
  /* TG68K_ALU.vhd:1268:17  */
  assign n11647 = div_bit ? n11645 : n11646;
  /* TG68K_ALU.vhd:1273:49  */
  assign n11648 = div_reg[30:0]; // extract
  /* TG68K_ALU.vhd:1273:63  */
  assign n11649 = ~div_bit;
  /* TG68K_ALU.vhd:1273:62  */
  assign n11650 = {n11648, n11649};
  /* TG68K_ALU.vhd:1276:66  */
  assign n11651 = div_quot[31:0]; // extract
  /* TG68K_ALU.vhd:1276:57  */
  assign n11653 = 32'b00000000000000000000000000000000 - n11651;
  /* TG68K_ALU.vhd:1279:64  */
  assign n11654 = div_quot[31:0]; // extract
  /* TG68K_ALU.vhd:1275:17  */
  assign n11655 = div_neg ? n11653 : n11654;
  /* TG68K_ALU.vhd:1282:44  */
  assign n11656 = ~div_bit;
  /* TG68K_ALU.vhd:1282:34  */
  assign n11657 = nozero | n11656;
  /* TG68K_ALU.vhd:1282:50  */
  assign n11658 = signedop & n11657;
  /* TG68K_ALU.vhd:1282:78  */
  assign n11659 = op2out[31]; // extract
  /* TG68K_ALU.vhd:1282:83  */
  assign n11660 = n11659 ^ op1_sign;
  /* TG68K_ALU.vhd:1282:96  */
  assign n11661 = n11660 ^ div_qsign;
  /* TG68K_ALU.vhd:1282:67  */
  assign n11662 = n11661 & n11658;
  /* TG68K_ALU.vhd:1283:37  */
  assign n11663 = ~signedop;
  /* TG68K_ALU.vhd:1283:54  */
  assign n11664 = div_over[32]; // extract
  /* TG68K_ALU.vhd:1283:58  */
  assign n11665 = ~n11664;
  /* TG68K_ALU.vhd:1283:42  */
  assign n11666 = n11665 & n11663;
  /* TG68K_ALU.vhd:1283:25  */
  assign n11667 = n11662 | n11666;
  /* TG68K_ALU.vhd:1283:65  */
  assign n11669 = 1'b1 & n11667;
  /* TG68K_ALU.vhd:1282:17  */
  assign n11672 = n11669 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1294:47  */
  assign n11678 = micro_state != 7'b1011010;
  /* TG68K_ALU.vhd:1298:47  */
  assign n11681 = micro_state == 7'b1010101;
  /* TG68K_ALU.vhd:1300:65  */
  assign n11682 = dividend[63]; // extract
  /* TG68K_ALU.vhd:1300:53  */
  assign n11683 = n11682 & divs;
  /* TG68K_ALU.vhd:1302:61  */
  assign n11685 = 64'b0000000000000000000000000000000000000000000000000000000000000000 - dividend;
  /* TG68K_ALU.vhd:1300:41  */
  assign n11686 = n11683 ? n11685 : dividend;
  /* TG68K_ALU.vhd:1300:41  */
  assign n11689 = n11683 ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1309:51  */
  assign n11690 = ~div_bit;
  /* TG68K_ALU.vhd:1309:63  */
  assign n11691 = n11690 | nozero;
  /* TG68K_ALU.vhd:1298:33  */
  assign n11692 = n11681 ? n11686 : div_quot;
  /* TG68K_ALU.vhd:1298:33  */
  assign n11694 = n11681 ? 1'b0 : n11691;
  /* TG68K_ALU.vhd:1311:47  */
  assign n11697 = micro_state == 7'b1010110;
  /* TG68K_ALU.vhd:1312:72  */
  assign n11698 = op2out[31]; // extract
  /* TG68K_ALU.vhd:1312:77  */
  assign n11699 = n11698 ^ op1_sign;
  /* TG68K_ALU.vhd:1312:61  */
  assign n11700 = signedop & n11699;
  /* TG68K_ALU.vhd:1316:73  */
  assign n11701 = div_reg[63:32]; // extract
  /* TG68K_ALU.vhd:1316:65  */
  assign n11703 = {1'b0, n11701};
  /* TG68K_ALU.vhd:1316:93  */
  assign n11705 = {1'b0, op2outext};
  /* TG68K_ALU.vhd:1316:123  */
  assign n11706 = op2out[15:0]; // extract
  /* TG68K_ALU.vhd:1316:116  */
  assign n11707 = {n11705, n11706};
  /* TG68K_ALU.vhd:1316:88  */
  assign n11708 = n11703 - n11707;
  /* TG68K_ALU.vhd:1319:40  */
  assign n11711 = exec[68]; // extract
  /* TG68K_ALU.vhd:1319:56  */
  assign n11712 = ~n11711;
  /* TG68K_ALU.vhd:1322:87  */
  assign n11713 = div_quot[63:32]; // extract
  /* TG68K_ALU.vhd:1322:78  */
  assign n11715 = 32'b00000000000000000000000000000000 - n11713;
  /* TG68K_ALU.vhd:1324:85  */
  assign n11716 = div_quot[63:32]; // extract
  /* TG68K_ALU.vhd:1321:41  */
  assign n11717 = op1_sign ? n11715 : n11716;
  assign n11718 = {n11717, result_div_pre};
  /* TG68K_ALU.vhd:1293:25  */
  assign n11720 = n11712 & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n11721 = n11678 & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n11723 = n11697 & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n11724 = n11697 & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n11727 = n11681 & clkena_lw;
  assign n11737 = {n9537, n9534};
  assign n11738 = {n9688, n9681, n9674};
  assign n11739 = {n9666, n9665, n9660, n9618};
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n11740 <= n11443;
  /* TG68K_ALU.vhd:996:17  */
  assign n11741 = {n9710, n9748};
  /* TG68K_ALU.vhd:1292:17  */
  assign n11742 = n11720 ? n11718 : result_div;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11743 <= n11742;
  /* TG68K_ALU.vhd:1292:17  */
  assign n11744 = n11721 ? n11672 : v_flag;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11745 <= n11744;
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n11746 <= n11444;
  /* TG68K_ALU.vhd:405:17  */
  assign n11748 = clkena_lw ? n9769 : bchg;
  /* TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n11749 <= n11748;
  /* TG68K_ALU.vhd:405:17  */
  assign n11750 = clkena_lw ? n9773 : bset;
  /* TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n11751 <= n11750;
  assign n11755 = mulu_reg[31:0]; // extract
  /* TG68K_ALU.vhd:1211:17  */
  assign n11756 = clkena_lw ? n11514 : n11755;
  /* TG68K_ALU.vhd:1211:17  */
  always @(posedge clk)
    n11757 <= n11756;
  assign n11759 = {32'bZ, n11757};
  /* TG68K_ALU.vhd:1292:17  */
  assign n11761 = clkena_lw ? n11692 : div_reg;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11762 <= n11761;
  /* TG68K_ALU.vhd:1292:17  */
  assign n11763 = {n11647, n11650};
  /* TG68K_ALU.vhd:1292:17  */
  assign n11765 = n11723 ? n11700 : div_neg;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11766 <= n11765;
  /* TG68K_ALU.vhd:1292:17  */
  assign n11767 = n11724 ? n11708 : div_over;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11768 <= n11767;
  /* TG68K_ALU.vhd:1292:17  */
  assign n11769 = clkena_lw ? n11694 : nozero;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11770 <= n11769;
  /* TG68K_ALU.vhd:1292:17  */
  assign n11771 = {n11623, n11620, n11618};
  /* TG68K_ALU.vhd:1292:17  */
  assign n11772 = clkena_lw ? divs : signedop;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11773 <= n11772;
  /* TG68K_ALU.vhd:1292:17  */
  assign n11774 = n11727 ? n11689 : op1_sign;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n11775 <= n11774;
  assign n11778 = {n10224, n10214, n10203, n10192, n10181, n10170, n10159, n10148, n10137, n10126, n10115, n10104, n10093, n10082, n10071, n10060, n10049, n10038, n10027, n10016, n10005, n9994, n9983, n9972, n9961, n9950, n9939, n9928, n9917, n9906, n9895, n9883};
  assign n11780 = {n10519, n10515, n10510, n10505, n10500, n10495, n10490, n10485, n10480, n10475, n10470, n10465, n10460, n10455, n10450, n10445, n10440, n10435, n10430, n10425, n10420, n10415, n10410, n10405, n10400, n10395, n10390, n10385, n10380, n10375, n10370, n10365, n10360, n10355, n10350, n10345, n10340, n10335, n10330, n10325};
  assign n11781 = {n10225, n10217, n10206, n10195, n10184, n10173, n10162, n10151, n10140, n10129, n10118, n10107, n10096, n10085, n10074, n10063, n10052, n10041, n10030, n10019, n10008, n9997, n9986, n9975, n9964, n9953, n9942, n9931, n9920, n9909, n9898, n9886};
  assign n11783 = {n10281, n10282};
  assign n11784 = {n10603, n10632, n10629};
  /* TG68K_ALU.vhd:446:17  */
  assign n11785 = clkena_lw ? n9832 : bf_bset;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11786 <= n11785;
  /* TG68K_ALU.vhd:446:17  */
  assign n11787 = clkena_lw ? n9836 : bf_bchg;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11788 <= n11787;
  /* TG68K_ALU.vhd:446:17  */
  assign n11789 = clkena_lw ? n9840 : bf_ins;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11790 <= n11789;
  /* TG68K_ALU.vhd:446:17  */
  assign n11791 = clkena_lw ? n9844 : bf_exts;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11792 <= n11791;
  /* TG68K_ALU.vhd:446:17  */
  assign n11793 = clkena_lw ? n9848 : bf_fffo;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11794 <= n11793;
  /* TG68K_ALU.vhd:446:17  */
  assign n11795 = clkena_lw ? n9857 : bf_d32;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11796 <= n11795;
  /* TG68K_ALU.vhd:446:17  */
  assign n11797 = clkena_lw ? n9851 : bf_s32;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11798 <= n11797;
  assign n11800 = {n11123, n11121, n11118, n11115, n11112, n11125};
  assign n11801 = {n10804, n10801, n10805, n10799, n10803};
  assign n11802 = {n11058, n11060};
  assign n11803 = {n11135, n11132, n11137};
  /* TG68K_ALU.vhd:446:17  */
  assign n11804 = clkena_lw ? n9859 : n11805;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n11805 <= n11804;
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n11806 <= n11447;
  /* TG68K_ALU.vhd:433:38  */
  assign n11807 = op1out[bit_number * 1 +: 1]; //(Bmux)
  /* TG68K_ALU.vhd:435:17  */
  assign n11808 = bit_number[4]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11809 = ~n11808;
  /* TG68K_ALU.vhd:435:17  */
  assign n11810 = bit_number[3]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11811 = ~n11810;
  /* TG68K_ALU.vhd:435:17  */
  assign n11812 = n11809 & n11811;
  /* TG68K_ALU.vhd:435:17  */
  assign n11813 = n11809 & n11810;
  /* TG68K_ALU.vhd:435:17  */
  assign n11814 = n11808 & n11811;
  /* TG68K_ALU.vhd:435:17  */
  assign n11815 = n11808 & n11810;
  /* TG68K_ALU.vhd:435:17  */
  assign n11816 = bit_number[2]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11817 = ~n11816;
  /* TG68K_ALU.vhd:435:17  */
  assign n11818 = n11812 & n11817;
  /* TG68K_ALU.vhd:435:17  */
  assign n11819 = n11812 & n11816;
  /* TG68K_ALU.vhd:435:17  */
  assign n11820 = n11813 & n11817;
  /* TG68K_ALU.vhd:435:17  */
  assign n11821 = n11813 & n11816;
  /* TG68K_ALU.vhd:435:17  */
  assign n11822 = n11814 & n11817;
  /* TG68K_ALU.vhd:435:17  */
  assign n11823 = n11814 & n11816;
  /* TG68K_ALU.vhd:435:17  */
  assign n11824 = n11815 & n11817;
  /* TG68K_ALU.vhd:435:17  */
  assign n11825 = n11815 & n11816;
  /* TG68K_ALU.vhd:435:17  */
  assign n11826 = bit_number[1]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11827 = ~n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11828 = n11818 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11829 = n11818 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11830 = n11819 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11831 = n11819 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11832 = n11820 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11833 = n11820 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11834 = n11821 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11835 = n11821 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11836 = n11822 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11837 = n11822 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11838 = n11823 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11839 = n11823 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11840 = n11824 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11841 = n11824 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11842 = n11825 & n11827;
  /* TG68K_ALU.vhd:435:17  */
  assign n11843 = n11825 & n11826;
  /* TG68K_ALU.vhd:435:17  */
  assign n11844 = bit_number[0]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11845 = ~n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11846 = n11828 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11847 = n11828 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11848 = n11829 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11849 = n11829 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11850 = n11830 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11851 = n11830 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11852 = n11831 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11853 = n11831 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11854 = n11832 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11855 = n11832 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11856 = n11833 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11857 = n11833 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11858 = n11834 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11859 = n11834 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11860 = n11835 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11861 = n11835 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11862 = n11836 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11863 = n11836 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11864 = n11837 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11865 = n11837 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11866 = n11838 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11867 = n11838 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11868 = n11839 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11869 = n11839 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11870 = n11840 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11871 = n11840 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11872 = n11841 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11873 = n11841 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11874 = n11842 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11875 = n11842 & n11844;
  /* TG68K_ALU.vhd:435:17  */
  assign n11876 = n11843 & n11845;
  /* TG68K_ALU.vhd:435:17  */
  assign n11877 = n11843 & n11844;
  /* TG68K_ALU.vhd:705:50  */
  assign n11878 = op1out[0]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11879 = n11846 ? n9805 : n11878;
  /* TG68K_ALU.vhd:705:41  */
  assign n11880 = op1out[1]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11881 = n11847 ? n9805 : n11880;
  /* TG68K_ALU.vhd:703:41  */
  assign n11882 = op1out[2]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11883 = n11848 ? n9805 : n11882;
  /* TG68K_ALU.vhd:702:48  */
  assign n11884 = op1out[3]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11885 = n11849 ? n9805 : n11884;
  /* TG68K_ALU.vhd:701:58  */
  assign n11886 = op1out[4]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11887 = n11850 ? n9805 : n11886;
  /* TG68K_ALU.vhd:695:50  */
  assign n11888 = op1out[5]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11889 = n11851 ? n9805 : n11888;
  assign n11890 = op1out[6]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11891 = n11852 ? n9805 : n11890;
  assign n11892 = op1out[7]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11893 = n11853 ? n9805 : n11892;
  assign n11894 = op1out[8]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11895 = n11854 ? n9805 : n11894;
  assign n11896 = op1out[9]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11897 = n11855 ? n9805 : n11896;
  /* TG68K_ALU.vhd:676:25  */
  assign n11898 = op1out[10]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11899 = n11856 ? n9805 : n11898;
  /* TG68K_ALU.vhd:678:65  */
  assign n11900 = op1out[11]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11901 = n11857 ? n9805 : n11900;
  /* TG68K_ALU.vhd:673:25  */
  assign n11902 = op1out[12]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11903 = n11858 ? n9805 : n11902;
  /* TG68K_ALU.vhd:670:25  */
  assign n11904 = op1out[13]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11905 = n11859 ? n9805 : n11904;
  /* TG68K_ALU.vhd:657:1  */
  assign n11906 = op1out[14]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11907 = n11860 ? n9805 : n11906;
  assign n11908 = op1out[15]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11909 = n11861 ? n9805 : n11908;
  assign n11910 = op1out[16]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11911 = n11862 ? n9805 : n11910;
  assign n11912 = op1out[17]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11913 = n11863 ? n9805 : n11912;
  assign n11914 = op1out[18]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11915 = n11864 ? n9805 : n11914;
  assign n11916 = op1out[19]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11917 = n11865 ? n9805 : n11916;
  assign n11918 = op1out[20]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11919 = n11866 ? n9805 : n11918;
  assign n11920 = op1out[21]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11921 = n11867 ? n9805 : n11920;
  assign n11922 = op1out[22]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11923 = n11868 ? n9805 : n11922;
  assign n11924 = op1out[23]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11925 = n11869 ? n9805 : n11924;
  assign n11926 = op1out[24]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11927 = n11870 ? n9805 : n11926;
  assign n11928 = op1out[25]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11929 = n11871 ? n9805 : n11928;
  assign n11930 = op1out[26]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11931 = n11872 ? n9805 : n11930;
  assign n11932 = op1out[27]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11933 = n11873 ? n9805 : n11932;
  assign n11934 = op1out[28]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11935 = n11874 ? n9805 : n11934;
  assign n11936 = op1out[29]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11937 = n11875 ? n9805 : n11936;
  assign n11938 = op1out[30]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11939 = n11876 ? n9805 : n11938;
  assign n11940 = op1out[31]; // extract
  /* TG68K_ALU.vhd:435:17  */
  assign n11941 = n11877 ? n9805 : n11940;
  assign n11942 = {n11941, n11939, n11937, n11935, n11933, n11931, n11929, n11927, n11925, n11923, n11921, n11919, n11917, n11915, n11913, n11911, n11909, n11907, n11905, n11903, n11901, n11899, n11897, n11895, n11893, n11891, n11889, n11887, n11885, n11883, n11881, n11879};
  /* TG68K_ALU.vhd:496:37  */
  assign n11943 = datareg[n10227 * 1 +: 1]; //(Bmux)
  /* TG68K_ALU.vhd:761:17  */
  assign n11944 = bit_msb[5]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n11945 = ~n11944;
  /* TG68K_ALU.vhd:761:17  */
  assign n11946 = bit_msb[4]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n11947 = ~n11946;
  /* TG68K_ALU.vhd:761:17  */
  assign n11948 = n11945 & n11947;
  /* TG68K_ALU.vhd:761:17  */
  assign n11949 = n11945 & n11946;
  /* TG68K_ALU.vhd:761:17  */
  assign n11950 = n11944 & n11947;
  /* TG68K_ALU.vhd:761:17  */
  assign n11951 = bit_msb[3]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n11952 = ~n11951;
  /* TG68K_ALU.vhd:761:17  */
  assign n11953 = n11948 & n11952;
  /* TG68K_ALU.vhd:761:17  */
  assign n11954 = n11948 & n11951;
  /* TG68K_ALU.vhd:761:17  */
  assign n11955 = n11949 & n11952;
  /* TG68K_ALU.vhd:761:17  */
  assign n11956 = n11949 & n11951;
  /* TG68K_ALU.vhd:761:17  */
  assign n11957 = n11950 & n11952;
  /* TG68K_ALU.vhd:761:17  */
  assign n11958 = bit_msb[2]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n11959 = ~n11958;
  /* TG68K_ALU.vhd:761:17  */
  assign n11960 = n11953 & n11959;
  /* TG68K_ALU.vhd:761:17  */
  assign n11961 = n11953 & n11958;
  /* TG68K_ALU.vhd:761:17  */
  assign n11962 = n11954 & n11959;
  /* TG68K_ALU.vhd:761:17  */
  assign n11963 = n11954 & n11958;
  /* TG68K_ALU.vhd:761:17  */
  assign n11964 = n11955 & n11959;
  /* TG68K_ALU.vhd:761:17  */
  assign n11965 = n11955 & n11958;
  /* TG68K_ALU.vhd:761:17  */
  assign n11966 = n11956 & n11959;
  /* TG68K_ALU.vhd:761:17  */
  assign n11967 = n11956 & n11958;
  /* TG68K_ALU.vhd:761:17  */
  assign n11968 = n11957 & n11959;
  /* TG68K_ALU.vhd:761:17  */
  assign n11969 = bit_msb[1]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n11970 = ~n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11971 = n11960 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11972 = n11960 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11973 = n11961 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11974 = n11961 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11975 = n11962 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11976 = n11962 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11977 = n11963 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11978 = n11963 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11979 = n11964 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11980 = n11964 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11981 = n11965 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11982 = n11965 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11983 = n11966 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11984 = n11966 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11985 = n11967 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11986 = n11967 & n11969;
  /* TG68K_ALU.vhd:761:17  */
  assign n11987 = n11968 & n11970;
  /* TG68K_ALU.vhd:761:17  */
  assign n11988 = bit_msb[0]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n11989 = ~n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n11990 = n11971 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n11991 = n11971 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n11992 = n11972 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n11993 = n11972 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n11994 = n11973 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n11995 = n11973 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n11996 = n11974 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n11997 = n11974 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n11998 = n11975 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n11999 = n11975 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12000 = n11976 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12001 = n11976 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12002 = n11977 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12003 = n11977 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12004 = n11978 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12005 = n11978 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12006 = n11979 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12007 = n11979 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12008 = n11980 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12009 = n11980 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12010 = n11981 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12011 = n11981 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12012 = n11982 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12013 = n11982 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12014 = n11983 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12015 = n11983 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12016 = n11984 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12017 = n11984 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12018 = n11985 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12019 = n11985 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12020 = n11986 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12021 = n11986 & n11988;
  /* TG68K_ALU.vhd:761:17  */
  assign n12022 = n11987 & n11989;
  /* TG68K_ALU.vhd:761:17  */
  assign n12023 = n11987 & n11988;
  assign n12024 = n10770[0]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12025 = n11990 ? 1'b1 : n12024;
  assign n12026 = n10770[1]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12027 = n11991 ? 1'b1 : n12026;
  assign n12028 = n10770[2]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12029 = n11992 ? 1'b1 : n12028;
  assign n12030 = n10770[3]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12031 = n11993 ? 1'b1 : n12030;
  /* TG68K_ALU.vhd:433:38  */
  assign n12032 = n10770[4]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12033 = n11994 ? 1'b1 : n12032;
  /* TG68K_ALU.vhd:405:17  */
  assign n12034 = n10770[5]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12035 = n11995 ? 1'b1 : n12034;
  assign n12036 = n10770[6]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12037 = n11996 ? 1'b1 : n12036;
  assign n12038 = n10770[7]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12039 = n11997 ? 1'b1 : n12038;
  /* TG68K_ALU.vhd:366:1  */
  assign n12040 = n10770[8]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12041 = n11998 ? 1'b1 : n12040;
  assign n12042 = n10770[9]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12043 = n11999 ? 1'b1 : n12042;
  assign n12044 = n10770[10]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12045 = n12000 ? 1'b1 : n12044;
  /* TG68K_ALU.vhd:210:1  */
  assign n12046 = n10770[11]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12047 = n12001 ? 1'b1 : n12046;
  /* TG68K_ALU.vhd:157:16  */
  assign n12048 = n10770[12]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12049 = n12002 ? 1'b1 : n12048;
  /* TG68K_ALU.vhd:150:16  */
  assign n12050 = n10770[13]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12051 = n12003 ? 1'b1 : n12050;
  /* TG68K_ALU.vhd:136:16  */
  assign n12052 = n10770[14]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12053 = n12004 ? 1'b1 : n12052;
  /* TG68K_ALU.vhd:128:16  */
  assign n12054 = n10770[15]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12055 = n12005 ? 1'b1 : n12054;
  /* TG68K_ALU.vhd:126:16  */
  assign n12056 = n10770[16]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12057 = n12006 ? 1'b1 : n12056;
  /* TG68K_ALU.vhd:114:16  */
  assign n12058 = n10770[17]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12059 = n12007 ? 1'b1 : n12058;
  /* TG68K_ALU.vhd:996:17  */
  assign n12060 = n10770[18]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12061 = n12008 ? 1'b1 : n12060;
  assign n12062 = n10770[19]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12063 = n12009 ? 1'b1 : n12062;
  assign n12064 = n10770[20]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12065 = n12010 ? 1'b1 : n12064;
  assign n12066 = n10770[21]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12067 = n12011 ? 1'b1 : n12066;
  assign n12068 = n10770[22]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12069 = n12012 ? 1'b1 : n12068;
  assign n12070 = n10770[23]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12071 = n12013 ? 1'b1 : n12070;
  assign n12072 = n10770[24]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12073 = n12014 ? 1'b1 : n12072;
  assign n12074 = n10770[25]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12075 = n12015 ? 1'b1 : n12074;
  assign n12076 = n10770[26]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12077 = n12016 ? 1'b1 : n12076;
  assign n12078 = n10770[27]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12079 = n12017 ? 1'b1 : n12078;
  assign n12080 = n10770[28]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12081 = n12018 ? 1'b1 : n12080;
  assign n12082 = n10770[29]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12083 = n12019 ? 1'b1 : n12082;
  assign n12084 = n10770[30]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12085 = n12020 ? 1'b1 : n12084;
  assign n12086 = n10770[31]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12087 = n12021 ? 1'b1 : n12086;
  assign n12088 = n10770[32]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12089 = n12022 ? 1'b1 : n12088;
  assign n12090 = n10770[33]; // extract
  /* TG68K_ALU.vhd:761:17  */
  assign n12091 = n12023 ? 1'b1 : n12090;
  assign n12092 = {n12091, n12089, n12087, n12085, n12083, n12081, n12079, n12077, n12075, n12073, n12071, n12069, n12067, n12065, n12063, n12061, n12059, n12057, n12055, n12053, n12051, n12049, n12047, n12045, n12043, n12041, n12039, n12037, n12035, n12033, n12031, n12029, n12027, n12025};
endmodule

module TG68KdotC_Kernel
  (input  clk,
   input  nReset,
   input  clkena_in,
   input  [15:0] data_in,
   input  [2:0] IPL,
   input  IPL_autovector,
   input  berr,
   input  [1:0] CPU,
   output [31:0] addr_out,
   output [15:0] data_write,
   output nWr,
   output nUDS,
   output nLDS,
   output [1:0] busstate,
   output longword,
   output nResetOut,
   output [2:0] FC,
   output clr_berr,
   output skipFetch,
   output [31:0] regin_out,
   output [3:0] CACR_out,
   output [31:0] VBR_out);
  wire use_vbr_stackframe;
  wire [3:0] syncreset;
  wire reset;
  wire clkena_lw;
  wire [31:0] tg68_pc;
  wire [31:0] tmp_tg68_pc;
  wire [31:0] tg68_pc_add;
  wire [31:0] pc_dataa;
  wire [31:0] pc_datab;
  wire [31:0] memaddr;
  wire [1:0] state;
  wire [1:0] datatype;
  wire [1:0] set_datatype;
  wire [1:0] exe_datatype;
  wire [1:0] setstate;
  wire setaddrvalue;
  wire addrvalue;
  wire [15:0] opcode;
  wire [15:0] exe_opcode;
  wire [15:0] sndopc;
  wire [31:0] exe_pc;
  wire [31:0] last_opc_pc;
  wire [15:0] last_opc_read;
  wire [31:0] reg_qa;
  wire [31:0] reg_qb;
  wire wwrena;
  wire lwrena;
  wire bwrena;
  wire regwrena_now;
  wire [3:0] rf_dest_addr;
  wire [3:0] rf_source_addr;
  wire [3:0] rf_source_addrd;
  wire [31:0] regin;
  wire [3:0] rdindex_a;
  wire [3:0] rdindex_b;
  wire wr_areg;
  wire [31:0] addr;
  wire [31:0] memaddr_reg;
  wire [31:0] memaddr_delta;
  wire [31:0] memaddr_delta_rega;
  wire [31:0] memaddr_delta_regb;
  wire use_base;
  wire [31:0] ea_data;
  wire [31:0] op1out;
  wire [31:0] op2out;
  wire [15:0] op1outbrief;
  wire [31:0] aluout;
  wire [31:0] data_write_tmp;
  wire [31:0] data_write_muxin;
  wire [47:0] data_write_mux;
  wire nextpass;
  wire setnextpass;
  wire setdispbyte;
  wire setdisp;
  wire regdirectsource;
  wire [31:0] addsub_q;
  wire [31:0] briefdata;
  wire [2:0] c_out;
  wire [31:0] memaddr_a;
  wire tg68_pc_brw;
  wire tg68_pc_word;
  wire getbrief;
  wire [15:0] brief;
  wire data_is_source;
  wire store_in_tmp;
  wire write_back;
  wire exec_write_back;
  wire setstackaddr;
  wire writepc;
  wire writepcbig;
  wire set_writepcbig;
  wire writepcnext;
  wire setopcode;
  wire decodeopc;
  wire execopc;
  wire execopc_alu;
  wire setexecopc;
  wire endopc;
  wire setendopc;
  wire [7:0] flags;
  wire [7:0] flagssr;
  wire [7:0] srin;
  wire exec_direct;
  wire exec_tas;
  wire set_exec_tas;
  wire exe_condition;
  wire ea_only;
  wire source_areg;
  wire source_lowbits;
  wire source_ldrlbits;
  wire source_ldrmbits;
  wire source_2ndhbits;
  wire source_2ndmbits;
  wire source_2ndlbits;
  wire dest_areg;
  wire dest_ldrareg;
  wire dest_ldrhbits;
  wire dest_ldrlbits;
  wire dest_2ndhbits;
  wire dest_2ndlbits;
  wire dest_hbits;
  wire [1:0] rot_bits;
  wire [1:0] set_rot_bits;
  wire [5:0] rot_cnt;
  wire [5:0] set_rot_cnt;
  wire movem_actiond;
  wire [3:0] movem_regaddr;
  wire [3:0] movem_mux;
  wire movem_presub;
  wire movem_run;
  wire set_direct_data;
  wire use_direct_data;
  wire direct_data;
  wire set_v_flag;
  wire set_vectoraddr;
  wire writesr;
  wire trap_berr;
  wire trap_illegal;
  wire trap_addr_error;
  wire trap_priv;
  wire trap_trace;
  wire trap_1010;
  wire trap_1111;
  wire trap_trap;
  wire trap_trapv;
  wire trap_interrupt;
  wire trapmake;
  wire trapd;
  wire [7:0] trap_sr;
  wire make_trace;
  wire make_berr;
  wire usestackframe2;
  wire set_stop;
  wire stop;
  wire [31:0] trap_vector;
  wire [31:0] trap_vector_vbr;
  wire [31:0] usp;
  wire [2:0] ipl_nr;
  wire [2:0] ripl_nr;
  wire [7:0] ipl_vec;
  wire interrupt;
  wire setinterrupt;
  wire svmode;
  wire presvmode;
  wire suppress_base;
  wire set_suppress_base;
  wire set_z_error;
  wire z_error;
  wire ea_build_now;
  wire build_logical;
  wire build_bcd;
  wire [31:0] data_read;
  wire [7:0] bf_ext_in;
  wire [7:0] bf_ext_out;
  wire long_start;
  wire long_start_alu;
  wire non_aligned;
  wire check_aligned;
  wire long_done;
  wire [5:0] memmask;
  wire [5:0] set_memmask;
  wire [3:0] memread;
  wire [5:0] wbmemmask;
  wire [5:0] memmaskmux;
  wire oddout;
  wire set_oddout;
  wire pcbase;
  wire set_pcbase;
  wire [31:0] last_data_read;
  wire [31:0] last_data_in;
  wire [5:0] bf_offset;
  wire [5:0] bf_width;
  wire [5:0] bf_bhits;
  wire [5:0] bf_shift;
  wire [5:0] alu_width;
  wire [5:0] alu_bf_shift;
  wire [5:0] bf_loffset;
  wire [31:0] bf_full_offset;
  wire [31:0] alu_bf_ffo_offset;
  wire [5:0] alu_bf_loffset;
  wire [31:0] movec_data;
  wire [31:0] vbr;
  wire [3:0] cacr;
  wire [2:0] dfc;
  wire [2:0] sfc;
  wire [88:0] set;
  wire [88:0] set_exec;
  wire [88:0] exec;
  wire [6:0] micro_state;
  wire [6:0] next_micro_state;
  wire [15:0] n15;
  wire [15:0] n16;
  wire [7:0] alu_n17;
  wire [4:0] n18;
  wire alu_n19;
  wire [7:0] alu_n20;
  wire [2:0] alu_n21;
  wire [31:0] alu_n22;
  wire [31:0] alu_n23;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire [1:0] n44;
  wire n46;
  wire [1:0] n47;
  wire n49;
  wire n50;
  wire n53;
  wire n58;
  wire n59;
  wire n62;
  wire n63;
  wire n65;
  wire [5:0] n66;
  wire [4:0] n67;
  wire [5:0] n69;
  wire n70;
  wire n71;
  wire n73;
  wire n74;
  wire n75;
  wire n78;
  wire n79;
  wire n83;
  wire [2:0] n85;
  wire [3:0] n87;
  wire n88;
  wire n89;
  wire n99;
  wire n101;
  wire n103;
  wire n106;
  wire n111;
  wire n112;
  wire [15:0] n113;
  wire [31:0] n114;
  wire [23:0] n115;
  wire [7:0] n116;
  wire [31:0] n117;
  wire [31:0] n118;
  wire n119;
  wire [1:0] n120;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire [3:0] n142;
  wire [3:0] n143;
  wire [3:0] n144;
  wire [3:0] n145;
  wire [15:0] n146;
  wire [15:0] n147;
  wire [15:0] n148;
  wire [15:0] n149;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire [7:0] n156;
  wire [7:0] n157;
  wire [7:0] n158;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire [3:0] n189;
  wire [3:0] n190;
  wire [3:0] n191;
  wire [3:0] n192;
  wire [15:0] n193;
  wire [15:0] n194;
  wire [15:0] n195;
  wire [15:0] n196;
  wire [15:0] n197;
  wire [31:0] n198;
  wire [31:0] n199;
  wire [15:0] n200;
  wire [31:0] n201;
  wire n202;
  wire [31:0] n203;
  wire [31:0] n205;
  wire [31:0] n206;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n217;
  wire [31:0] n218;
  wire n219;
  wire n220;
  wire [15:0] n222;
  wire [47:0] n223;
  wire [39:0] n224;
  wire [47:0] n226;
  wire [47:0] n227;
  wire n228;
  wire n229;
  wire [15:0] n230;
  wire n231;
  wire n232;
  wire [15:0] n233;
  wire [1:0] n234;
  wire n236;
  wire [7:0] n237;
  wire [7:0] n238;
  wire [15:0] n239;
  wire [1:0] n240;
  wire n242;
  wire [7:0] n243;
  wire [7:0] n244;
  wire [15:0] n245;
  wire [15:0] n246;
  wire [15:0] n247;
  wire [15:0] n248;
  wire [15:0] n249;
  wire [15:0] n250;
  wire n251;
  wire [7:0] n252;
  wire [7:0] n253;
  wire [7:0] n254;
  wire [7:0] n255;
  wire n268;
  wire n276;
  wire n279;
  wire n283;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire [31:0] n298;
  wire [31:0] n299;
  wire [31:0] n300;
  wire [31:0] n301;
  wire [7:0] n302;
  wire [7:0] n303;
  wire [7:0] n304;
  wire [15:0] n305;
  wire [7:0] n306;
  wire n307;
  wire [15:0] n308;
  wire [15:0] n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n317;
  wire n318;
  wire n321;
  wire n323;
  wire [1:0] n324;
  reg n327;
  reg n330;
  wire n333;
  wire n335;
  wire n337;
  wire n339;
  wire n341;
  wire n343;
  wire n345;
  wire n348;
  wire n351;
  wire n356;
  wire n357;
  wire [3:0] n358;
  wire n359;
  wire [2:0] n360;
  wire [3:0] n362;
  wire [2:0] n363;
  wire [3:0] n364;
  wire [3:0] n365;
  wire [2:0] n366;
  wire [3:0] n368;
  wire [2:0] n369;
  wire [3:0] n371;
  wire [2:0] n372;
  wire [3:0] n373;
  wire [2:0] n374;
  wire n376;
  wire n377;
  wire [2:0] n378;
  wire [3:0] n379;
  wire [2:0] n380;
  wire [3:0] n382;
  wire [3:0] n383;
  wire [3:0] n384;
  wire [3:0] n386;
  wire [3:0] n387;
  wire [3:0] n388;
  wire [3:0] n389;
  wire [3:0] n390;
  wire [3:0] n391;
  wire [3:0] n392;
  wire [3:0] n393;
  wire n397;
  wire n398;
  wire n399;
  wire [3:0] n401;
  wire [3:0] n402;
  wire [2:0] n403;
  wire [3:0] n405;
  wire [2:0] n406;
  wire [3:0] n408;
  wire [2:0] n409;
  wire [3:0] n411;
  wire [2:0] n412;
  wire [3:0] n414;
  wire [2:0] n415;
  wire [3:0] n417;
  wire [2:0] n418;
  wire [3:0] n419;
  wire n420;
  wire [2:0] n421;
  wire [3:0] n422;
  wire [3:0] n424;
  wire [3:0] n425;
  wire [3:0] n426;
  wire [3:0] n427;
  wire [3:0] n428;
  wire [3:0] n429;
  wire [3:0] n430;
  wire [3:0] n431;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire [31:0] n444;
  wire [31:0] n445;
  wire [31:0] n447;
  wire [15:0] n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire [3:0] n468;
  wire [3:0] n469;
  wire [3:0] n470;
  wire [3:0] n471;
  wire [15:0] n472;
  wire n473;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire [7:0] n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire [3:0] n495;
  wire [3:0] n496;
  wire [7:0] n497;
  wire n498;
  wire [2:0] n499;
  wire [2:0] n500;
  wire n502;
  wire n505;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire [15:0] n512;
  wire [15:0] n513;
  wire [15:0] n514;
  wire [15:0] n515;
  wire [15:0] n516;
  wire [31:0] n517;
  wire [15:0] n518;
  wire [15:0] n519;
  wire [15:0] n520;
  wire [15:0] n521;
  wire [15:0] n522;
  wire [31:0] n523;
  wire [31:0] n524;
  wire [31:0] n525;
  wire [15:0] n526;
  wire [15:0] n527;
  wire [15:0] n528;
  wire [15:0] n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire [3:0] n555;
  wire [3:0] n556;
  wire [3:0] n557;
  wire [3:0] n558;
  wire [3:0] n559;
  wire [3:0] n560;
  wire [15:0] n561;
  wire [7:0] n562;
  wire [23:0] n563;
  wire [7:0] n564;
  wire [23:0] n565;
  wire [23:0] n566;
  wire [7:0] n567;
  wire n572;
  wire n574;
  wire n575;
  wire n576;
  wire n578;
  wire n580;
  wire n583;
  wire n585;
  wire n587;
  wire n588;
  wire n590;
  wire n591;
  wire n593;
  wire n595;
  wire n596;
  wire n597;
  wire n599;
  wire n601;
  wire n602;
  wire n604;
  wire n606;
  wire n608;
  wire n609;
  wire n611;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n620;
  wire n621;
  wire n622;
  wire [31:0] n623;
  wire [31:0] n624;
  wire [31:0] n625;
  wire n626;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n634;
  wire [11:0] n635;
  wire [15:0] n637;
  wire [11:0] n638;
  wire [15:0] n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire [15:0] n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n652;
  wire n653;
  wire n654;
  wire [23:0] n655;
  wire [23:0] n656;
  wire [23:0] n657;
  wire [7:0] n658;
  wire n659;
  wire [15:0] n660;
  wire [15:0] n661;
  wire [15:0] n662;
  wire [15:0] n663;
  wire [15:0] n664;
  wire [15:0] n665;
  wire [15:0] n666;
  wire [31:0] n667;
  wire [31:0] n668;
  wire [15:0] n669;
  wire [15:0] n670;
  wire [15:0] n671;
  wire [15:0] n672;
  wire [15:0] n673;
  wire [31:0] n674;
  wire [31:0] n675;
  wire [31:0] n676;
  wire [31:0] n677;
  wire [31:0] n678;
  wire [31:0] n679;
  wire [31:0] n680;
  wire [15:0] n681;
  wire [15:0] n682;
  wire [15:0] n683;
  wire [15:0] n684;
  wire [15:0] n685;
  wire n686;
  wire [31:0] n687;
  wire [31:0] n688;
  wire n689;
  wire n692;
  wire [31:0] n693;
  wire n694;
  wire n696;
  wire [31:0] n697;
  wire n698;
  wire n700;
  wire [31:0] n702;
  wire [31:0] n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire [31:0] n711;
  wire [31:0] n712;
  wire n714;
  wire n716;
  wire n717;
  wire n719;
  wire n721;
  wire n722;
  wire n724;
  wire n737;
  wire [15:0] n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire [3:0] n755;
  wire [3:0] n756;
  wire [3:0] n757;
  wire [3:0] n758;
  wire [15:0] n759;
  wire [15:0] n760;
  wire [15:0] n761;
  wire [31:0] n762;
  wire n763;
  wire n765;
  wire n767;
  wire [1:0] n768;
  wire [15:0] n769;
  wire [31:0] n770;
  wire n772;
  wire [14:0] n773;
  wire [15:0] n774;
  wire [30:0] n775;
  wire [31:0] n777;
  wire n779;
  wire [13:0] n780;
  wire [15:0] n781;
  wire [29:0] n782;
  wire [31:0] n784;
  wire n786;
  wire [12:0] n787;
  wire [15:0] n788;
  wire [28:0] n789;
  wire [31:0] n791;
  wire n793;
  wire [3:0] n794;
  reg [31:0] n795;
  wire [31:0] n796;
  wire [9:0] n803;
  wire [9:0] n804;
  wire [9:0] n806;
  wire [9:0] n808;
  wire [9:0] n810;
  wire n811;
  wire [9:0] n813;
  wire [9:0] n815;
  wire [9:0] n817;
  wire [9:0] n819;
  wire [9:0] n821;
  wire [9:0] n823;
  wire [3:0] n824;
  wire [7:0] n826;
  wire [9:0] n828;
  wire [9:0] n829;
  wire n830;
  wire [9:0] n832;
  wire [9:0] n833;
  wire [31:0] n834;
  wire [31:0] n837;
  wire [31:0] n838;
  wire n840;
  wire n841;
  wire n842;
  wire [2:0] n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire [3:0] n852;
  wire [3:0] n853;
  wire [7:0] n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire [3:0] n871;
  wire [3:0] n872;
  wire [3:0] n873;
  wire [3:0] n874;
  wire [15:0] n875;
  wire n876;
  wire [31:0] n877;
  wire [7:0] n878;
  wire [7:0] n879;
  wire [7:0] n880;
  wire [23:0] n881;
  wire [23:0] n882;
  wire [23:0] n883;
  wire [31:0] n884;
  wire [31:0] n885;
  wire n886;
  wire n887;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire [4:0] n896;
  wire [4:0] n897;
  wire [3:0] n899;
  wire [4:0] n901;
  wire [4:0] n902;
  wire [4:0] n903;
  wire [4:0] n904;
  wire [4:0] n905;
  wire [26:0] n906;
  wire [26:0] n907;
  wire [26:0] n908;
  wire n910;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n925;
  wire n926;
  wire n927;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n936;
  wire [31:0] n937;
  wire n939;
  wire [31:0] n940;
  wire [31:0] n942;
  wire n944;
  wire [31:0] n945;
  wire [31:0] n947;
  wire n949;
  wire [31:0] n950;
  wire [31:0] n952;
  wire n954;
  wire [31:0] n955;
  wire [31:0] n957;
  wire n959;
  wire [31:0] n960;
  wire [31:0] n962;
  wire n964;
  wire [31:0] n965;
  wire [31:0] n967;
  wire n969;
  wire [31:0] n970;
  wire [31:0] n972;
  wire n975;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n983;
  wire n984;
  wire [31:0] n993;
  wire [31:0] n994;
  wire [31:0] n995;
  wire n996;
  wire [31:0] n998;
  wire [31:0] n1002;
  localparam [2:0] n1003 = 3'b000;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire [3:0] n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire [3:0] n1018;
  wire [3:0] n1019;
  wire [7:0] n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire [3:0] n1037;
  wire [3:0] n1038;
  wire [3:0] n1039;
  wire [3:0] n1040;
  wire [15:0] n1041;
  wire [1:0] n1043;
  wire [1:0] n1044;
  wire n1045;
  wire n1046;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1063;
  wire n1065;
  wire n1067;
  wire n1068;
  wire [2:0] n1069;
  wire n1070;
  wire n1071;
  wire [1:0] n1072;
  wire n1073;
  wire [1:0] n1074;
  wire [1:0] n1075;
  wire [7:0] n1077;
  wire [7:0] n1078;
  wire [7:0] n1079;
  wire [23:0] n1080;
  wire [23:0] n1081;
  wire [23:0] n1082;
  wire [31:0] n1083;
  wire [31:0] n1084;
  wire [31:0] n1085;
  wire [31:0] n1086;
  wire n1088;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire [2:0] n1105;
  wire n1106;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1115;
  wire n1117;
  wire n1120;
  wire n1122;
  wire n1126;
  wire n1129;
  wire n1132;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1147;
  wire [2:0] n1149;
  wire [3:0] n1151;
  wire [5:0] n1153;
  wire [1:0] n1154;
  wire [1:0] n1155;
  wire [3:0] n1156;
  wire n1157;
  wire n1158;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire [31:0] n1164;
  wire [31:0] n1165;
  wire [31:0] n1166;
  wire [31:0] n1167;
  wire [5:0] n1168;
  wire [3:0] n1169;
  wire n1170;
  wire n1171;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire [7:0] n1178;
  wire n1181;
  wire n1184;
  wire [2:0] n1185;
  wire [7:0] n1186;
  wire n1188;
  wire n1192;
  wire n1195;
  wire [2:0] n1197;
  wire [7:0] n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1203;
  wire [2:0] n1204;
  wire [7:0] n1205;
  wire n1207;
  wire n1208;
  wire n1209;
  wire [7:0] n1210;
  wire [7:0] n1211;
  wire n1213;
  wire [15:0] n1214;
  wire [31:0] n1215;
  wire [15:0] n1216;
  wire [7:0] n1217;
  wire n1219;
  wire [7:0] n1220;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1226;
  wire n1228;
  wire n1230;
  wire n1232;
  wire n1234;
  wire n1235;
  wire [31:0] n1236;
  wire [31:0] n1237;
  wire [31:0] n1239;
  wire [5:0] n1240;
  wire [5:0] n1241;
  wire [31:0] n1242;
  wire [5:0] n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire [1:0] n1256;
  wire [1:0] n1257;
  wire n1259;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1266;
  wire n1268;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1275;
  wire n1276;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1298;
  wire [5:0] n1301;
  wire [5:0] n1304;
  wire n1306;
  wire [5:0] n1308;
  wire [5:0] n1310;
  wire n1312;
  wire [5:0] n1313;
  wire [5:0] n1314;
  wire n1315;
  wire [5:0] n1317;
  wire [5:0] n1319;
  wire n1320;
  wire [1:0] n1321;
  wire [1:0] n1323;
  wire n1325;
  wire [5:0] n1326;
  wire [5:0] n1327;
  wire n1328;
  wire [1:0] n1329;
  wire [1:0] n1331;
  wire n1333;
  wire [5:0] n1335;
  wire [5:0] n1336;
  wire n1337;
  wire n1338;
  wire n1340;
  wire [1:0] n1341;
  wire n1342;
  wire n1343;
  wire n1345;
  wire n1346;
  wire [5:0] n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1353;
  wire n1355;
  wire n1356;
  wire [15:0] n1357;
  wire [15:0] n1358;
  wire [15:0] n1359;
  wire n1360;
  wire n1361;
  wire n1363;
  wire [15:0] n1364;
  wire [15:0] n1365;
  wire [31:0] n1366;
  wire n1367;
  wire n1368;
  wire n1370;
  wire [15:0] n1372;
  wire n1374;
  wire [15:0] n1375;
  wire [31:0] n1376;
  wire n1378;
  wire n1379;
  wire [7:0] n1380;
  wire [1:0] n1381;
  wire [1:0] n1382;
  wire [1:0] n1383;
  wire [1:0] n1384;
  wire n1385;
  wire [15:0] n1386;
  wire [15:0] n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire [7:0] n1408;
  wire n1409;
  wire n1410;
  wire [5:0] n1411;
  wire [3:0] n1413;
  wire [5:0] n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire [1:0] n1420;
  wire [1:0] n1421;
  wire [31:0] n1423;
  wire [1:0] n1425;
  wire [1:0] n1426;
  wire n1428;
  wire [15:0] n1430;
  wire [15:0] n1431;
  wire [31:0] n1432;
  wire [31:0] n1433;
  wire [15:0] n1435;
  wire n1436;
  wire n1438;
  wire [15:0] n1439;
  wire n1441;
  wire n1443;
  wire n1445;
  wire n1447;
  wire n1449;
  wire [1:0] n1450;
  wire [5:0] n1452;
  wire n1454;
  wire n1456;
  wire n1458;
  wire [7:0] n1459;
  wire n1461;
  wire n1463;
  wire [2:0] n1464;
  wire [7:0] n1465;
  wire n1467;
  wire n1469;
  wire [5:0] n1471;
  wire [3:0] n1472;
  wire [5:0] n1473;
  wire n1474;
  wire [5:0] n1475;
  wire [5:0] n1476;
  wire [31:0] n1477;
  wire [5:0] n1478;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1525;
  wire n1526;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1534;
  wire n1535;
  wire n1536;
  wire [1:0] n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire [35:0] n1541;
  wire [47:0] n1542;
  wire [88:0] n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire [84:0] n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire [1:0] n1556;
  wire n1558;
  wire [88:0] n1560;
  wire [88:0] n1561;
  wire [88:0] n1562;
  wire n1563;
  wire n1564;
  wire [16:0] n1565;
  wire [70:0] n1566;
  wire [88:0] n1568;
  wire n1576;
  wire [4:0] n1577;
  wire [5:0] n1579;
  wire [4:0] n1580;
  wire [5:0] n1582;
  wire [5:0] n1583;
  wire n1584;
  wire [4:0] n1585;
  localparam [31:0] n1586 = 32'b00000000000000000000000000000000;
  wire [26:0] n1587;
  wire [31:0] n1588;
  wire [31:0] n1589;
  wire n1591;
  wire [4:0] n1592;
  wire [4:0] n1594;
  wire [4:0] n1595;
  wire [4:0] n1597;
  wire [4:0] n1598;
  wire [5:0] n1599;
  wire n1600;
  wire n1601;
  wire [2:0] n1602;
  wire n1604;
  wire [5:0] n1606;
  wire [5:0] n1607;
  wire [4:0] n1609;
  wire [1:0] n1610;
  wire n1612;
  wire [2:0] n1613;
  wire n1615;
  wire [5:0] n1617;
  wire [5:0] n1619;
  wire [5:0] n1620;
  wire [4:0] n1622;
  wire [2:0] n1623;
  wire n1625;
  wire [2:0] n1626;
  wire [5:0] n1628;
  wire [5:0] n1630;
  wire [4:0] n1632;
  wire [2:0] n1633;
  wire [2:0] n1635;
  wire [5:0] n1637;
  wire [5:0] n1638;
  wire [5:0] n1639;
  wire [1:0] n1641;
  wire [1:0] n1642;
  wire n1643;
  wire [2:0] n1644;
  wire [5:0] n1645;
  wire [5:0] n1646;
  wire [2:0] n1647;
  wire n1649;
  wire n1651;
  wire n1653;
  wire n1655;
  wire [3:0] n1656;
  reg [5:0] n1662;
  wire n1664;
  wire [5:0] n1666;
  wire n1670;
  wire [7:0] n1671;
  wire [7:0] n1672;
  wire n1673;
  wire [7:0] n1674;
  wire [7:0] n1675;
  wire n1676;
  wire [7:0] n1677;
  wire [7:0] n1678;
  wire [7:0] n1679;
  wire [7:0] n1680;
  wire [7:0] n1681;
  wire [7:0] n1682;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1697;
  wire n1698;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1711;
  wire n1713;
  wire n1715;
  wire n1716;
  wire n1718;
  wire n1719;
  wire n1720;
  wire [7:0] n1721;
  wire [4:0] n1722;
  wire n1723;
  wire [7:0] n1724;
  wire [7:0] n1725;
  wire n1726;
  wire [2:0] n1727;
  wire [2:0] n1728;
  wire [4:0] n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire [7:0] n1736;
  wire [7:0] n1737;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1750;
  wire n1751;
  wire [2:0] n1753;
  wire n1754;
  wire n1755;
  wire [7:0] n1756;
  wire [7:0] n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire [7:0] n1763;
  wire n1765;
  wire n1767;
  wire n1769;
  wire [1:0] n1779;
  wire n1781;
  wire [5:0] n1783;
  wire [5:0] n1785;
  localparam [88:0] n1788 = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [1:0] n1791;
  wire n1793;
  wire n1795;
  wire [1:0] n1796;
  reg [1:0] n1800;
  wire n1801;
  wire n1803;
  wire n1804;
  wire n1807;
  wire n1808;
  wire n1810;
  wire n1811;
  wire [1:0] n1814;
  wire n1817;
  wire [6:0] n1822;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire [6:0] n1833;
  wire n1834;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1840;
  wire [1:0] n1842;
  wire n1844;
  wire n1845;
  wire [6:0] n1848;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire [6:0] n1857;
  wire n1858;
  wire n1860;
  wire [1:0] n1862;
  wire n1863;
  wire [6:0] n1864;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1871;
  wire [1:0] n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1879;
  wire n1880;
  wire [1:0] n1883;
  wire n1884;
  wire [6:0] n1886;
  wire n1887;
  wire n1892;
  wire [1:0] n1894;
  wire [1:0] n1895;
  wire [1:0] n1896;
  wire n1899;
  wire n1900;
  wire n1901;
  wire [1:0] n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1908;
  wire n1909;
  wire n1912;
  wire n1913;
  wire n1914;
  wire [2:0] n1915;
  wire n1917;
  wire [2:0] n1919;
  wire n1921;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1928;
  wire n1929;
  wire [2:0] n1931;
  wire n1933;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1940;
  wire n1942;
  wire n1943;
  wire n1945;
  wire n1946;
  wire n1948;
  wire n1950;
  wire [2:0] n1951;
  wire n1953;
  wire n1956;
  wire n1959;
  wire n1962;
  wire n1964;
  wire n1966;
  wire n1968;
  wire [4:0] n1969;
  reg n1972;
  reg n1975;
  reg n1978;
  reg n1982;
  reg n1986;
  wire n1987;
  reg n1988;
  reg n1989;
  reg [6:0] n1994;
  wire n1996;
  wire [3:0] n1997;
  reg n2000;
  reg n2003;
  reg n2005;
  reg n2007;
  reg n2009;
  wire n2010;
  reg n2011;
  wire n2012;
  reg n2013;
  wire n2014;
  reg n2015;
  wire n2016;
  reg n2017;
  wire n2018;
  reg n2019;
  reg n2020;
  reg [6:0] n2023;
  wire n2025;
  wire n2028;
  wire n2031;
  wire n2034;
  wire n2037;
  wire [1:0] n2039;
  wire n2040;
  wire n2041;
  wire [1:0] n2042;
  wire [1:0] n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire [1:0] n2054;
  wire [1:0] n2055;
  wire [6:0] n2057;
  wire [3:0] n2058;
  wire n2059;
  wire [2:0] n2060;
  wire n2062;
  wire n2063;
  wire n2066;
  wire n2067;
  wire n2071;
  wire n2072;
  wire n2074;
  wire n2076;
  wire n2077;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2083;
  wire n2084;
  wire n2085;
  wire [6:0] n2087;
  wire n2090;
  wire n2091;
  wire [2:0] n2092;
  wire n2094;
  wire n2095;
  wire [2:0] n2096;
  wire n2098;
  wire [5:0] n2099;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire [6:0] n2106;
  wire n2108;
  wire [1:0] n2109;
  wire n2111;
  wire n2112;
  wire n2113;
  wire [1:0] n2114;
  wire n2116;
  wire [2:0] n2117;
  wire n2119;
  wire n2120;
  wire [1:0] n2121;
  wire n2123;
  wire n2124;
  wire n2125;
  wire [1:0] n2128;
  wire n2130;
  wire [1:0] n2131;
  wire n2133;
  wire n2136;
  wire n2139;
  wire n2141;
  wire [1:0] n2142;
  wire n2144;
  wire [1:0] n2147;
  wire n2148;
  wire n2149;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire [6:0] n2157;
  wire n2160;
  wire n2162;
  wire n2164;
  wire n2165;
  wire [1:0] n2166;
  wire n2168;
  wire n2171;
  wire n2174;
  wire n2176;
  wire n2178;
  wire n2180;
  wire n2182;
  wire n2184;
  wire n2186;
  wire n2187;
  wire [2:0] n2188;
  wire n2190;
  wire n2191;
  wire n2192;
  wire [1:0] n2193;
  wire n2195;
  wire [1:0] n2196;
  wire n2198;
  wire n2199;
  wire [2:0] n2200;
  wire n2202;
  wire [1:0] n2203;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire [5:0] n2209;
  wire n2211;
  wire n2212;
  wire n2213;
  wire [1:0] n2214;
  wire n2216;
  wire n2218;
  wire [1:0] n2219;
  reg [1:0] n2223;
  wire n2224;
  wire [5:0] n2225;
  wire n2227;
  wire n2228;
  wire n2230;
  wire n2231;
  wire [6:0] n2233;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire [6:0] n2241;
  wire n2243;
  wire n2244;
  wire [1:0] n2250;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire [6:0] n2263;
  wire [1:0] n2264;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire [6:0] n2278;
  wire [1:0] n2279;
  wire [1:0] n2280;
  wire n2282;
  wire n2285;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire [6:0] n2301;
  wire [1:0] n2302;
  wire n2304;
  wire [1:0] n2305;
  wire n2307;
  wire n2308;
  wire [2:0] n2309;
  wire n2311;
  wire n2312;
  wire [2:0] n2313;
  wire n2315;
  wire n2316;
  wire [3:0] n2317;
  wire n2319;
  wire n2320;
  wire [1:0] n2322;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire [6:0] n2330;
  wire n2331;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2339;
  wire n2340;
  wire n2343;
  wire n2346;
  wire [1:0] n2348;
  wire n2350;
  wire n2351;
  wire n2352;
  wire [6:0] n2354;
  wire [1:0] n2355;
  wire n2356;
  wire n2359;
  wire n2362;
  wire n2364;
  wire [1:0] n2365;
  wire n2367;
  wire [1:0] n2368;
  wire [1:0] n2369;
  wire n2371;
  wire n2373;
  wire n2375;
  wire [6:0] n2376;
  wire [1:0] n2377;
  wire [1:0] n2378;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2384;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2402;
  wire n2404;
  wire [6:0] n2405;
  wire [1:0] n2406;
  wire [1:0] n2407;
  wire n2409;
  wire n2411;
  wire n2413;
  wire n2415;
  wire [1:0] n2416;
  wire [1:0] n2417;
  wire n2419;
  wire n2420;
  wire n2421;
  wire [1:0] n2422;
  wire [1:0] n2423;
  wire [1:0] n2424;
  wire [1:0] n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2431;
  wire n2433;
  wire [6:0] n2434;
  wire [2:0] n2435;
  wire n2437;
  wire n2438;
  wire [1:0] n2439;
  wire n2441;
  wire n2442;
  wire [1:0] n2443;
  wire n2445;
  wire n2446;
  wire [2:0] n2447;
  wire n2449;
  wire [1:0] n2450;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2457;
  wire n2460;
  wire n2462;
  wire n2464;
  wire [1:0] n2465;
  wire n2467;
  wire [2:0] n2468;
  wire n2470;
  wire n2471;
  wire [2:0] n2472;
  wire n2474;
  wire [2:0] n2475;
  wire n2477;
  wire [1:0] n2478;
  wire n2480;
  wire n2481;
  wire [2:0] n2482;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2492;
  wire n2495;
  wire n2497;
  wire n2499;
  wire n2501;
  wire n2503;
  wire [2:0] n2504;
  wire n2506;
  wire [2:0] n2507;
  wire n2509;
  wire [1:0] n2510;
  wire n2512;
  wire n2513;
  wire [2:0] n2514;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2523;
  wire n2525;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2531;
  wire [2:0] n2532;
  wire n2534;
  wire [2:0] n2535;
  wire n2537;
  wire n2538;
  wire [2:0] n2539;
  wire n2541;
  wire [1:0] n2542;
  wire n2544;
  wire n2545;
  wire n2548;
  wire n2550;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2556;
  wire [2:0] n2557;
  wire n2559;
  wire [2:0] n2560;
  wire n2562;
  wire [1:0] n2563;
  wire n2565;
  wire n2566;
  wire [2:0] n2567;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2576;
  wire n2578;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2584;
  wire [2:0] n2585;
  wire n2587;
  wire [2:0] n2588;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2596;
  wire n2598;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire [5:0] n2616;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2631;
  wire n2633;
  wire n2634;
  wire n2636;
  wire n2637;
  wire n2638;
  wire [1:0] n2640;
  wire [2:0] n2641;
  wire [1:0] n2642;
  wire [2:0] n2643;
  wire [2:0] n2644;
  wire [1:0] n2645;
  wire [1:0] n2646;
  wire [6:0] n2648;
  wire [1:0] n2649;
  wire n2652;
  wire n2654;
  wire [2:0] n2655;
  wire [2:0] n2656;
  wire n2657;
  wire n2658;
  wire [1:0] n2659;
  wire [1:0] n2660;
  wire [6:0] n2661;
  wire n2662;
  wire n2663;
  wire [5:0] n2664;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2678;
  wire n2680;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire [6:0] n2689;
  wire [1:0] n2690;
  wire n2692;
  wire n2695;
  wire [2:0] n2696;
  wire n2698;
  wire [1:0] n2699;
  wire n2701;
  wire n2704;
  wire n2707;
  wire n2709;
  wire [1:0] n2710;
  wire n2712;
  wire n2714;
  wire n2715;
  wire n2717;
  wire n2718;
  wire n2720;
  wire n2722;
  wire n2724;
  wire n2726;
  wire n2728;
  wire n2729;
  wire n2731;
  wire n2733;
  wire n2734;
  wire [1:0] n2735;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2741;
  wire n2742;
  wire [2:0] n2743;
  wire [2:0] n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire [1:0] n2749;
  wire [1:0] n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2757;
  wire n2759;
  wire [6:0] n2760;
  wire n2761;
  wire n2763;
  wire n2764;
  wire n2766;
  wire n2768;
  wire n2770;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2776;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2785;
  wire n2787;
  wire [6:0] n2788;
  wire n2789;
  wire n2791;
  wire n2792;
  wire n2794;
  wire n2796;
  wire n2798;
  wire n2800;
  wire n2802;
  wire n2804;
  wire n2806;
  wire n2808;
  wire n2810;
  wire n2811;
  wire [3:0] n2812;
  wire n2814;
  wire [3:0] n2816;
  wire n2818;
  wire n2820;
  wire n2821;
  wire [1:0] n2822;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2829;
  wire [2:0] n2830;
  wire [2:0] n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire [1:0] n2836;
  wire [1:0] n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2844;
  wire [3:0] n2846;
  wire n2848;
  wire n2850;
  wire [6:0] n2851;
  wire n2852;
  wire [1:0] n2853;
  wire n2855;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2861;
  wire n2862;
  wire n2864;
  wire [2:0] n2865;
  wire [2:0] n2866;
  wire n2868;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire [1:0] n2878;
  wire [1:0] n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2888;
  wire n2890;
  wire n2892;
  wire n2894;
  wire [3:0] n2896;
  wire n2898;
  wire n2900;
  wire [6:0] n2901;
  wire [1:0] n2902;
  wire [1:0] n2903;
  wire n2904;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2910;
  wire n2911;
  wire n2913;
  wire n2915;
  wire [1:0] n2916;
  wire [1:0] n2917;
  wire [2:0] n2918;
  wire [2:0] n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire [1:0] n2931;
  wire [1:0] n2932;
  wire [1:0] n2933;
  wire [1:0] n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2944;
  wire [3:0] n2946;
  wire n2948;
  wire n2949;
  wire n2950;
  wire [6:0] n2951;
  wire [1:0] n2953;
  wire [1:0] n2954;
  wire n2956;
  wire n2958;
  wire n2960;
  wire n2961;
  wire n2963;
  wire n2965;
  wire n2967;
  wire n2969;
  wire n2971;
  wire [1:0] n2972;
  wire [1:0] n2973;
  wire [2:0] n2974;
  wire [2:0] n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire [1:0] n2982;
  wire [1:0] n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire [1:0] n2988;
  wire [1:0] n2989;
  wire [1:0] n2990;
  wire [1:0] n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3002;
  wire n3004;
  wire [3:0] n3006;
  wire n3008;
  wire n3010;
  wire n3011;
  wire [6:0] n3012;
  wire n3014;
  wire [1:0] n3015;
  wire n3017;
  wire [2:0] n3018;
  wire n3020;
  wire n3021;
  wire [3:0] n3022;
  wire n3024;
  wire [1:0] n3025;
  wire n3027;
  wire n3028;
  wire n3029;
  wire n3030;
  wire [2:0] n3031;
  wire n3033;
  wire [2:0] n3034;
  wire n3036;
  wire n3037;
  wire n3038;
  wire n3039;
  wire [2:0] n3041;
  wire n3043;
  wire n3045;
  wire n3046;
  wire [1:0] n3047;
  wire n3049;
  wire [1:0] n3050;
  wire n3052;
  wire n3055;
  wire n3057;
  wire [1:0] n3058;
  wire n3060;
  wire n3062;
  wire [1:0] n3063;
  reg [1:0] n3067;
  wire n3068;
  wire n3071;
  wire [1:0] n3072;
  wire n3074;
  wire n3075;
  wire [2:0] n3076;
  wire n3078;
  wire n3081;
  wire n3083;
  wire n3086;
  wire n3088;
  wire [1:0] n3089;
  wire n3091;
  wire n3092;
  wire n3093;
  wire n3094;
  wire [2:0] n3095;
  wire n3098;
  wire n3100;
  wire n3101;
  wire n3102;
  wire [2:0] n3104;
  wire n3106;
  wire n3108;
  wire n3109;
  wire n3110;
  wire n3111;
  wire n3112;
  wire [2:0] n3114;
  wire n3116;
  wire n3118;
  wire n3119;
  wire n3120;
  wire n3121;
  wire n3122;
  wire n3124;
  wire n3125;
  wire n3127;
  wire n3129;
  wire n3130;
  wire n3132;
  wire n3133;
  wire n3135;
  wire n3137;
  wire [2:0] n3138;
  wire n3140;
  wire n3143;
  wire [1:0] n3144;
  reg n3145;
  reg [6:0] n3148;
  wire n3150;
  wire [4:0] n3151;
  reg [1:0] n3153;
  reg n3155;
  wire n3156;
  reg n3157;
  wire n3158;
  reg n3159;
  wire n3160;
  reg n3161;
  reg n3162;
  reg n3163;
  reg n3164;
  reg [6:0] n3168;
  wire [1:0] n3169;
  wire n3170;
  wire [1:0] n3171;
  wire n3172;
  wire n3173;
  wire [1:0] n3174;
  wire n3175;
  wire n3176;
  wire n3177;
  wire [6:0] n3178;
  wire [1:0] n3179;
  wire n3180;
  wire n3181;
  wire n3183;
  wire n3186;
  wire n3188;
  wire n3190;
  wire n3193;
  wire n3196;
  wire n3199;
  wire [1:0] n3200;
  wire n3202;
  wire n3203;
  wire n3204;
  wire [1:0] n3205;
  wire [1:0] n3206;
  wire n3207;
  wire n3209;
  wire n3211;
  wire n3212;
  wire n3214;
  wire n3216;
  wire n3217;
  wire n3219;
  wire n3220;
  wire n3221;
  wire n3222;
  wire [2:0] n3223;
  wire n3225;
  wire [2:0] n3226;
  wire n3228;
  wire n3229;
  wire n3230;
  wire n3231;
  wire n3232;
  wire n3239;
  wire n3242;
  wire n3245;
  wire n3247;
  wire n3249;
  wire n3251;
  wire n3253;
  wire n3254;
  wire n3255;
  wire [1:0] n3256;
  wire n3258;
  wire n3259;
  wire n3260;
  wire [2:0] n3261;
  wire n3263;
  wire n3264;
  wire [3:0] n3265;
  wire n3267;
  wire n3268;
  wire [2:0] n3272;
  wire n3274;
  wire n3277;
  wire n3280;
  wire n3283;
  wire n3284;
  wire [1:0] n3286;
  wire n3288;
  wire n3290;
  wire n3292;
  wire n3293;
  wire n3296;
  wire n3299;
  wire n3302;
  wire n3304;
  wire n3306;
  wire n3307;
  wire n3310;
  wire n3313;
  wire n3315;
  wire n3316;
  wire n3317;
  wire n3319;
  wire n3321;
  wire [1:0] n3322;
  wire n3324;
  wire n3326;
  wire n3327;
  wire n3329;
  wire n3331;
  wire n3332;
  wire n3333;
  wire n3334;
  wire n3336;
  wire n3337;
  wire n3338;
  wire n3339;
  wire n3341;
  wire n3342;
  wire n3344;
  wire [2:0] n3345;
  wire n3347;
  wire [3:0] n3348;
  wire n3350;
  wire [1:0] n3351;
  wire n3353;
  wire n3354;
  wire n3355;
  wire n3356;
  wire n3358;
  wire n3359;
  wire n3360;
  wire n3361;
  wire n3362;
  wire n3363;
  wire n3364;
  wire n3365;
  wire n3368;
  wire n3369;
  wire n3371;
  wire n3372;
  wire n3373;
  wire n3374;
  wire n3375;
  wire n3376;
  wire n3377;
  wire n3378;
  wire n3381;
  wire [1:0] n3383;
  wire n3386;
  wire n3388;
  wire n3389;
  wire n3390;
  wire [1:0] n3392;
  wire n3394;
  wire n3395;
  wire n3396;
  wire n3397;
  wire n3398;
  wire n3399;
  wire [1:0] n3400;
  wire n3402;
  wire n3403;
  wire n3404;
  wire n3405;
  wire n3406;
  wire n3408;
  wire n3409;
  wire n3412;
  wire n3416;
  wire n3419;
  wire n3421;
  wire n3423;
  wire n3426;
  wire n3427;
  wire n3428;
  wire n3430;
  wire [1:0] n3431;
  wire n3433;
  wire n3435;
  wire n3437;
  wire n3439;
  wire n3441;
  wire n3442;
  wire n3443;
  wire n3445;
  wire n3447;
  wire [1:0] n3448;
  wire [1:0] n3449;
  wire n3451;
  wire n3453;
  wire n3454;
  wire n3456;
  wire n3457;
  wire n3458;
  wire n3459;
  wire n3460;
  wire n3461;
  wire n3462;
  wire n3463;
  wire n3464;
  wire n3465;
  wire n3466;
  wire n3467;
  wire n3469;
  wire n3471;
  wire n3473;
  wire n3475;
  wire n3477;
  wire [2:0] n3478;
  wire [2:0] n3479;
  wire n3481;
  wire [2:0] n3482;
  wire n3484;
  wire [1:0] n3485;
  wire n3487;
  wire n3488;
  wire n3489;
  wire [1:0] n3490;
  wire n3492;
  wire n3493;
  wire n3494;
  wire n3496;
  wire n3498;
  wire n3499;
  wire n3501;
  wire n3503;
  wire n3504;
  wire n3505;
  wire n3506;
  wire n3508;
  wire [1:0] n3509;
  wire n3511;
  wire n3514;
  wire n3515;
  wire [1:0] n3517;
  wire n3520;
  wire n3523;
  wire n3526;
  wire n3529;
  wire n3531;
  wire n3533;
  wire [1:0] n3537;
  wire n3539;
  wire n3542;
  wire n3544;
  wire n3545;
  wire n3546;
  wire n3547;
  wire n3549;
  wire n3552;
  wire n3554;
  wire n3556;
  wire n3558;
  wire n3559;
  wire n3560;
  wire n3561;
  wire n3562;
  wire n3564;
  wire n3566;
  wire n3568;
  wire n3569;
  wire n3570;
  wire n3571;
  wire n3573;
  wire n3575;
  wire n3578;
  wire n3580;
  wire n3582;
  wire n3584;
  wire n3585;
  wire n3586;
  wire n3587;
  wire n3588;
  wire [1:0] n3589;
  wire [1:0] n3591;
  wire n3593;
  wire n3595;
  wire n3597;
  wire [2:0] n3598;
  wire n3600;
  wire [2:0] n3601;
  wire n3603;
  wire [1:0] n3604;
  wire n3606;
  wire n3607;
  wire n3608;
  wire [1:0] n3609;
  wire n3611;
  wire n3612;
  wire n3614;
  wire n3616;
  wire [1:0] n3618;
  wire n3620;
  wire n3623;
  wire [1:0] n3625;
  wire n3628;
  wire n3631;
  wire n3634;
  wire n3637;
  wire n3639;
  wire n3641;
  wire n3643;
  wire n3645;
  wire n3646;
  wire n3647;
  wire n3648;
  wire n3650;
  wire n3652;
  wire n3653;
  wire [1:0] n3654;
  wire n3656;
  wire n3659;
  wire n3660;
  wire n3661;
  wire n3663;
  wire n3665;
  wire n3667;
  wire n3669;
  wire n3670;
  wire n3671;
  wire n3673;
  wire n3675;
  wire n3676;
  wire n3677;
  wire n3678;
  wire n3680;
  wire n3682;
  wire n3684;
  wire n3686;
  wire n3687;
  wire n3688;
  wire n3690;
  wire n3692;
  wire n3694;
  wire n3696;
  wire [1:0] n3697;
  wire n3699;
  wire [2:0] n3700;
  wire n3702;
  wire [3:0] n3703;
  wire n3705;
  wire [1:0] n3706;
  wire n3708;
  wire n3709;
  wire n3710;
  wire [1:0] n3711;
  wire n3713;
  wire n3714;
  wire n3716;
  wire n3717;
  wire n3718;
  wire n3719;
  wire n3720;
  wire n3722;
  wire n3723;
  wire [1:0] n3725;
  wire n3728;
  wire n3731;
  wire n3734;
  wire n3737;
  wire n3739;
  wire [2:0] n3740;
  wire n3742;
  wire [2:0] n3743;
  wire n3745;
  wire [1:0] n3746;
  wire n3748;
  wire n3749;
  wire n3750;
  wire [1:0] n3753;
  wire n3755;
  wire n3758;
  wire n3760;
  wire n3761;
  wire n3764;
  wire n3767;
  wire n3770;
  wire n3773;
  wire n3776;
  wire n3778;
  wire n3779;
  wire n3780;
  wire n3782;
  wire n3784;
  wire n3785;
  wire n3787;
  wire n3788;
  wire n3789;
  wire n3790;
  wire n3791;
  wire n3793;
  wire n3794;
  wire n3795;
  wire n3796;
  wire n3797;
  wire n3799;
  wire n3801;
  wire n3803;
  wire [1:0] n3804;
  wire n3806;
  wire [2:0] n3807;
  wire n3809;
  wire [3:0] n3810;
  wire n3812;
  wire [1:0] n3813;
  wire n3815;
  wire n3816;
  wire n3817;
  wire [1:0] n3818;
  wire n3820;
  wire n3821;
  wire n3823;
  wire n3824;
  wire n3825;
  wire n3826;
  wire n3827;
  wire [1:0] n3830;
  wire [1:0] n3831;
  wire [1:0] n3832;
  wire n3833;
  wire [1:0] n3834;
  wire n3836;
  wire n3837;
  wire n3838;
  wire n3840;
  wire n3841;
  wire n3842;
  wire n3843;
  wire n3844;
  wire [1:0] n3846;
  wire [1:0] n3848;
  wire n3849;
  wire n3852;
  wire n3855;
  wire n3858;
  wire n3861;
  wire n3863;
  wire n3864;
  wire n3865;
  wire n3867;
  wire n3870;
  wire n3872;
  wire n3874;
  wire n3876;
  wire n3878;
  wire [2:0] n3879;
  wire n3881;
  wire [2:0] n3882;
  wire n3884;
  wire [1:0] n3885;
  wire n3887;
  wire n3888;
  wire n3889;
  wire [2:0] n3892;
  wire n3894;
  wire n3897;
  wire n3899;
  wire n3900;
  wire n3903;
  wire n3906;
  wire n3909;
  wire n3912;
  wire n3914;
  wire n3916;
  wire n3918;
  wire n3920;
  wire n3921;
  wire n3922;
  wire n3924;
  wire n3926;
  wire n3927;
  wire n3929;
  wire n3930;
  wire n3931;
  wire n3933;
  wire n3934;
  wire n3935;
  wire n3937;
  wire n3939;
  wire n3941;
  wire n3943;
  wire n3944;
  wire [2:0] n3945;
  wire n3947;
  wire n3948;
  wire n3949;
  wire n3950;
  wire n3954;
  wire n3955;
  wire [1:0] n3958;
  wire n3960;
  wire n3961;
  wire n3962;
  wire [1:0] n3963;
  wire n3965;
  wire n3966;
  wire [2:0] n3967;
  wire n3969;
  wire [1:0] n3970;
  wire n3972;
  wire n3973;
  wire n3974;
  wire n3975;
  wire n3976;
  wire n3977;
  wire [1:0] n3978;
  wire n3980;
  wire [2:0] n3981;
  wire n3983;
  wire n3984;
  wire [3:0] n3985;
  wire n3987;
  wire n3988;
  wire n3989;
  wire n3990;
  wire n3992;
  wire n3993;
  wire [1:0] n3995;
  wire [2:0] n3996;
  wire n3998;
  wire [2:0] n3999;
  wire n4001;
  wire n4002;
  wire n4004;
  wire n4005;
  wire n4009;
  wire n4011;
  wire [2:0] n4012;
  wire n4014;
  wire n4018;
  wire n4019;
  wire n4020;
  wire n4022;
  wire n4023;
  wire n4024;
  wire n4027;
  wire n4028;
  wire n4029;
  wire n4030;
  wire [2:0] n4032;
  wire n4034;
  wire [2:0] n4035;
  wire n4037;
  wire n4038;
  wire [2:0] n4039;
  wire n4041;
  wire n4042;
  wire n4044;
  wire n4045;
  wire [6:0] n4048;
  wire n4049;
  wire n4050;
  wire n4051;
  wire n4052;
  wire [6:0] n4053;
  wire n4054;
  wire n4056;
  wire n4057;
  wire [1:0] n4061;
  wire n4062;
  wire n4063;
  wire [1:0] n4066;
  wire n4068;
  wire n4069;
  wire n4070;
  wire n4071;
  wire n4072;
  wire [6:0] n4074;
  wire [1:0] n4075;
  wire n4077;
  wire n4079;
  wire n4081;
  wire n4082;
  wire n4083;
  wire n4084;
  wire n4087;
  wire n4089;
  wire n4092;
  wire n4095;
  wire [1:0] n4096;
  wire n4098;
  wire n4100;
  wire n4102;
  wire n4104;
  wire [1:0] n4105;
  wire n4107;
  wire n4109;
  wire n4111;
  wire n4113;
  wire n4115;
  wire [6:0] n4116;
  wire [1:0] n4117;
  wire [1:0] n4118;
  wire n4120;
  wire n4123;
  wire n4125;
  wire n4127;
  wire n4129;
  wire n4130;
  wire n4131;
  wire n4132;
  wire n4133;
  wire n4134;
  wire n4135;
  wire n4136;
  wire n4137;
  wire [1:0] n4138;
  wire n4139;
  wire n4140;
  wire n4141;
  wire n4142;
  wire n4143;
  wire n4144;
  wire n4146;
  wire n4148;
  wire n4150;
  wire n4151;
  wire n4153;
  wire [6:0] n4154;
  wire n4155;
  wire [1:0] n4156;
  wire n4158;
  wire [2:0] n4159;
  wire n4161;
  wire n4162;
  wire [3:0] n4163;
  wire n4165;
  wire [1:0] n4166;
  wire n4168;
  wire n4169;
  wire n4170;
  wire n4172;
  wire n4173;
  wire n4174;
  wire n4175;
  wire n4177;
  wire n4179;
  wire n4180;
  wire n4181;
  wire n4184;
  wire n4185;
  wire n4186;
  wire n4187;
  wire [6:0] n4189;
  wire n4191;
  wire n4192;
  wire [1:0] n4193;
  wire n4195;
  wire n4196;
  wire n4197;
  wire n4198;
  wire n4201;
  wire [1:0] n4203;
  wire [6:0] n4205;
  wire n4209;
  wire n4212;
  wire n4213;
  wire n4214;
  wire n4215;
  wire n4216;
  wire n4217;
  wire n4218;
  wire n4219;
  wire [1:0] n4220;
  wire n4222;
  wire [2:0] n4223;
  wire n4225;
  wire n4226;
  wire [3:0] n4227;
  wire n4229;
  wire [1:0] n4230;
  wire n4232;
  wire n4233;
  wire n4234;
  wire n4235;
  wire n4236;
  wire n4238;
  wire n4240;
  wire n4241;
  wire n4242;
  wire n4243;
  wire n4244;
  wire n4246;
  wire n4248;
  wire n4249;
  wire n4250;
  wire n4251;
  wire n4254;
  wire n4255;
  wire n4256;
  wire n4257;
  wire [6:0] n4259;
  wire n4261;
  wire n4262;
  wire [1:0] n4263;
  wire n4265;
  wire n4266;
  wire n4267;
  wire n4268;
  wire n4269;
  wire n4271;
  wire n4272;
  wire [6:0] n4275;
  wire [1:0] n4277;
  wire n4280;
  wire n4283;
  wire n4284;
  wire n4285;
  wire [6:0] n4286;
  wire [1:0] n4287;
  wire n4289;
  wire n4290;
  wire n4291;
  wire n4294;
  wire [1:0] n4296;
  wire n4297;
  wire n4300;
  wire n4302;
  wire n4304;
  wire n4306;
  wire n4309;
  wire n4312;
  wire n4314;
  wire n4316;
  wire n4318;
  wire [6:0] n4319;
  wire [1:0] n4321;
  wire [1:0] n4322;
  wire n4324;
  wire n4326;
  wire n4327;
  wire n4329;
  wire n4331;
  wire n4333;
  wire n4335;
  wire n4336;
  wire n4337;
  wire n4339;
  wire n4340;
  wire n4342;
  wire n4343;
  wire [6:0] n4344;
  wire n4345;
  wire [2:0] n4346;
  wire n4348;
  wire [2:0] n4351;
  wire n4353;
  wire n4354;
  wire [1:0] n4355;
  wire n4357;
  wire n4358;
  wire [2:0] n4359;
  wire n4361;
  wire n4362;
  wire [3:0] n4363;
  wire n4365;
  wire n4366;
  wire n4368;
  wire n4369;
  wire [1:0] n4372;
  wire n4374;
  wire n4375;
  wire n4376;
  wire [6:0] n4378;
  wire n4379;
  wire [1:0] n4381;
  wire [1:0] n4382;
  wire n4383;
  wire n4386;
  wire n4389;
  wire n4392;
  wire n4395;
  wire n4397;
  wire n4398;
  wire [1:0] n4399;
  wire n4400;
  wire n4402;
  wire n4404;
  wire n4406;
  wire n4408;
  wire n4409;
  wire n4410;
  wire [6:0] n4411;
  wire [1:0] n4412;
  wire n4413;
  wire n4415;
  wire n4417;
  wire n4419;
  wire n4421;
  wire n4422;
  wire n4423;
  wire n4425;
  wire n4427;
  wire [6:0] n4428;
  wire [2:0] n4429;
  wire n4431;
  wire n4441;
  wire n4444;
  wire n4447;
  wire n4448;
  wire n4449;
  wire n4450;
  wire n4451;
  wire n4452;
  wire n4453;
  wire n4454;
  wire n4455;
  wire n4456;
  wire [6:0] n4458;
  wire [2:0] n4459;
  wire n4461;
  wire [2:0] n4462;
  wire n4464;
  wire [1:0] n4465;
  wire n4467;
  wire n4468;
  wire n4469;
  wire [1:0] n4474;
  wire n4476;
  wire n4479;
  wire n4481;
  wire n4482;
  wire n4485;
  wire n4488;
  wire n4491;
  wire n4494;
  wire n4497;
  wire n4499;
  wire n4500;
  wire n4501;
  wire n4503;
  wire n4505;
  wire n4507;
  wire n4509;
  wire [1:0] n4511;
  wire n4513;
  wire n4514;
  wire n4516;
  wire n4517;
  wire n4519;
  wire n4521;
  wire n4523;
  wire n4525;
  wire n4527;
  wire n4529;
  wire n4530;
  wire n4531;
  wire n4532;
  wire n4533;
  wire n4535;
  wire n4536;
  wire n4537;
  wire n4538;
  wire n4539;
  wire n4541;
  wire n4543;
  wire n4544;
  wire n4545;
  wire [1:0] n4547;
  wire [1:0] n4548;
  wire n4550;
  wire n4551;
  wire n4553;
  wire n4555;
  wire n4557;
  wire n4558;
  wire n4559;
  wire n4560;
  wire [2:0] n4561;
  wire n4562;
  wire n4563;
  wire n4564;
  wire n4565;
  wire n4566;
  wire n4567;
  wire n4568;
  wire [2:0] n4569;
  wire [2:0] n4570;
  wire n4571;
  wire n4573;
  wire n4575;
  wire n4577;
  wire n4579;
  wire n4580;
  wire [6:0] n4581;
  wire [1:0] n4582;
  wire [1:0] n4583;
  wire n4585;
  wire n4586;
  wire n4588;
  wire n4590;
  wire n4591;
  wire n4593;
  wire n4595;
  wire n4597;
  wire n4598;
  wire n4599;
  wire n4601;
  wire n4603;
  wire n4604;
  wire n4605;
  wire n4607;
  wire n4608;
  wire n4609;
  wire n4610;
  wire n4611;
  wire n4612;
  wire n4613;
  wire n4614;
  wire n4615;
  wire n4616;
  wire n4617;
  wire [2:0] n4618;
  wire [2:0] n4619;
  wire n4621;
  wire n4622;
  wire n4623;
  wire n4624;
  wire n4626;
  wire n4628;
  wire n4630;
  wire n4632;
  wire n4634;
  wire [6:0] n4635;
  wire [1:0] n4636;
  wire [1:0] n4637;
  wire n4639;
  wire n4640;
  wire n4641;
  wire n4643;
  wire n4644;
  wire n4646;
  wire n4648;
  wire n4650;
  wire n4652;
  wire n4653;
  wire n4654;
  wire n4656;
  wire n4657;
  wire n4658;
  wire n4659;
  wire n4660;
  wire n4661;
  wire n4662;
  wire n4663;
  wire n4664;
  wire n4665;
  wire n4666;
  wire n4667;
  wire n4668;
  wire n4669;
  wire n4670;
  wire n4671;
  wire n4672;
  wire n4673;
  wire n4674;
  wire n4675;
  wire n4676;
  wire n4677;
  wire n4678;
  wire n4679;
  wire n4680;
  wire n4681;
  wire n4682;
  wire n4683;
  wire n4684;
  wire n4685;
  wire n4686;
  wire n4687;
  wire n4688;
  wire n4689;
  wire n4690;
  wire n4691;
  wire n4693;
  wire n4695;
  wire n4697;
  wire n4699;
  wire n4701;
  wire n4703;
  wire n4705;
  wire n4706;
  wire n4708;
  wire [6:0] n4709;
  wire n4711;
  wire n4713;
  wire n4714;
  wire [4:0] n4715;
  wire n4717;
  wire [1:0] n4718;
  wire n4720;
  wire n4721;
  wire [1:0] n4722;
  wire n4724;
  wire [2:0] n4725;
  wire n4727;
  wire [2:0] n4728;
  wire n4730;
  wire [1:0] n4731;
  wire n4733;
  wire n4734;
  wire n4735;
  wire n4736;
  wire [1:0] n4737;
  wire n4739;
  wire [2:0] n4740;
  wire n4742;
  wire n4743;
  wire [3:0] n4744;
  wire n4746;
  wire [1:0] n4747;
  wire n4749;
  wire n4750;
  wire n4751;
  wire n4752;
  wire n4753;
  wire n4756;
  wire n4758;
  wire n4761;
  wire [1:0] n4763;
  wire n4765;
  wire [1:0] n4766;
  wire n4768;
  wire n4771;
  wire [1:0] n4773;
  wire n4776;
  wire n4779;
  wire n4781;
  wire n4782;
  wire n4784;
  wire n4786;
  wire n4788;
  wire n4790;
  wire n4793;
  wire n4796;
  wire n4799;
  wire n4801;
  wire n4803;
  wire [1:0] n4804;
  wire n4806;
  wire n4808;
  wire n4810;
  wire n4812;
  wire n4814;
  wire n4816;
  wire n4818;
  wire n4820;
  wire n4822;
  wire n4824;
  wire n4825;
  wire n4826;
  wire [1:0] n4827;
  wire n4829;
  wire n4830;
  wire [2:0] n4831;
  wire n4833;
  wire n4834;
  wire [3:0] n4835;
  wire n4837;
  wire n4838;
  wire n4839;
  wire [6:0] n4841;
  wire n4843;
  wire n4844;
  wire n4845;
  wire n4846;
  wire n4847;
  wire [1:0] n4850;
  wire n4852;
  wire n4853;
  wire n4854;
  wire [6:0] n4856;
  wire n4858;
  wire n4859;
  wire n4860;
  wire n4861;
  wire n4863;
  wire n4865;
  wire n4868;
  wire n4870;
  wire n4871;
  wire n4872;
  wire n4873;
  wire n4875;
  wire n4877;
  wire [1:0] n4879;
  wire n4880;
  wire n4881;
  wire n4882;
  wire [1:0] n4884;
  wire [1:0] n4885;
  wire n4886;
  wire n4888;
  wire n4891;
  wire n4894;
  wire n4897;
  wire n4900;
  wire [1:0] n4901;
  wire n4903;
  wire [1:0] n4904;
  wire [6:0] n4905;
  wire [6:0] n4906;
  wire n4908;
  wire n4910;
  wire n4911;
  wire n4913;
  wire n4914;
  wire n4916;
  wire n4917;
  wire n4919;
  wire n4920;
  wire n4922;
  wire n4923;
  wire n4925;
  wire n4926;
  wire n4928;
  wire n4929;
  wire n4931;
  wire n4932;
  wire n4934;
  wire n4935;
  wire n4937;
  wire n4938;
  wire n4940;
  wire n4941;
  wire n4943;
  wire n4944;
  wire n4946;
  wire n4947;
  wire n4949;
  wire n4950;
  wire n4952;
  wire n4953;
  wire n4961;
  wire n4964;
  wire n4967;
  wire n4968;
  wire n4969;
  wire n4970;
  wire n4971;
  wire n4972;
  wire n4973;
  wire [6:0] n4975;
  wire n4977;
  wire n4979;
  wire n4980;
  wire n4982;
  wire n4983;
  wire n4985;
  wire n4986;
  wire n4988;
  wire n4989;
  wire n4991;
  wire n4992;
  wire n4994;
  wire n4995;
  wire n4997;
  wire n4998;
  wire [1:0] n5005;
  wire n5007;
  wire n5010;
  wire n5013;
  wire n5014;
  wire n5015;
  wire n5016;
  wire n5017;
  wire [6:0] n5019;
  wire n5021;
  wire n5023;
  wire n5024;
  wire n5026;
  wire n5027;
  wire n5029;
  wire n5030;
  wire n5032;
  wire n5033;
  wire n5035;
  wire n5036;
  wire n5038;
  wire n5039;
  wire n5041;
  wire n5042;
  wire [1:0] n5045;
  wire n5048;
  wire n5051;
  wire n5054;
  wire n5057;
  wire n5058;
  wire n5059;
  wire n5061;
  wire n5063;
  wire n5064;
  wire n5066;
  wire n5067;
  wire n5069;
  wire n5070;
  wire n5072;
  wire n5073;
  wire n5075;
  wire n5076;
  wire n5078;
  wire n5079;
  wire n5081;
  wire n5082;
  wire [1:0] n5086;
  wire n5089;
  wire n5092;
  wire n5093;
  wire n5094;
  wire n5096;
  wire n5098;
  wire n5100;
  wire n5101;
  wire n5103;
  wire n5104;
  wire n5106;
  wire n5107;
  wire n5109;
  wire n5110;
  wire n5112;
  wire n5113;
  wire n5115;
  wire n5116;
  wire n5118;
  wire n5119;
  wire n5120;
  wire [5:0] n5124;
  wire n5125;
  wire n5126;
  wire [5:0] n5127;
  wire n5130;
  wire n5133;
  wire n5134;
  wire n5135;
  wire n5136;
  wire n5137;
  wire n5139;
  wire n5141;
  wire n5142;
  wire n5144;
  wire n5147;
  wire n5149;
  wire n5150;
  wire n5151;
  wire n5154;
  wire n5157;
  wire n5159;
  wire n5161;
  wire n5162;
  wire n5163;
  wire n5165;
  wire n5168;
  wire n5169;
  wire n5170;
  wire n5171;
  wire [1:0] n5173;
  wire n5175;
  wire [1:0] n5176;
  wire n5177;
  wire n5178;
  wire [1:0] n5179;
  wire [1:0] n5180;
  wire [6:0] n5182;
  wire n5183;
  wire n5184;
  wire n5187;
  wire n5190;
  wire n5192;
  wire n5194;
  wire n5195;
  wire n5197;
  wire n5199;
  wire n5200;
  wire [1:0] n5205;
  wire n5207;
  wire n5209;
  wire [1:0] n5210;
  wire n5211;
  wire n5212;
  wire [1:0] n5213;
  wire [1:0] n5214;
  wire [6:0] n5216;
  wire n5218;
  wire [1:0] n5223;
  wire n5225;
  wire [1:0] n5226;
  wire n5227;
  wire n5228;
  wire [1:0] n5229;
  wire [1:0] n5230;
  wire [6:0] n5232;
  wire n5234;
  wire [1:0] n5236;
  wire n5237;
  wire n5239;
  wire n5240;
  wire n5243;
  wire n5246;
  wire n5248;
  wire n5250;
  wire n5251;
  wire [11:0] n5252;
  wire n5254;
  wire n5256;
  wire n5258;
  wire n5259;
  wire [1:0] n5260;
  wire [1:0] n5261;
  wire n5262;
  wire n5263;
  wire n5267;
  wire n5269;
  wire n5271;
  wire [6:0] n5273;
  wire [1:0] n5275;
  wire n5276;
  wire n5279;
  wire n5282;
  wire [1:0] n5283;
  wire [1:0] n5284;
  wire [1:0] n5286;
  wire [6:0] n5287;
  wire [1:0] n5288;
  wire n5289;
  wire n5292;
  wire n5294;
  wire n5296;
  wire [1:0] n5297;
  wire [1:0] n5299;
  wire [6:0] n5300;
  wire n5302;
  wire n5304;
  wire n5305;
  wire [12:0] n5306;
  reg n5307;
  reg [1:0] n5312;
  reg [1:0] n5313;
  reg n5314;
  reg n5315;
  reg n5316;
  reg n5318;
  reg n5320;
  reg [5:0] n5321;
  reg n5322;
  reg n5325;
  reg n5327;
  reg n5330;
  reg n5332;
  reg n5336;
  reg n5338;
  wire n5339;
  reg n5340;
  wire n5341;
  reg n5342;
  wire n5343;
  reg n5344;
  wire n5345;
  reg n5346;
  wire n5347;
  reg n5348;
  wire n5349;
  reg n5350;
  wire n5351;
  reg n5352;
  wire n5353;
  reg n5354;
  wire [1:0] n5355;
  reg [1:0] n5356;
  wire [1:0] n5357;
  reg [1:0] n5358;
  wire n5359;
  wire n5360;
  reg n5361;
  wire n5362;
  wire n5363;
  reg n5364;
  wire n5365;
  reg n5366;
  reg n5368;
  reg n5370;
  reg [1:0] n5372;
  reg n5374;
  reg [6:0] n5375;
  wire n5376;
  wire [1:0] n5377;
  wire [1:0] n5378;
  wire n5379;
  wire n5380;
  wire n5381;
  wire n5383;
  wire n5385;
  wire n5387;
  wire n5389;
  wire [5:0] n5390;
  wire n5391;
  wire n5392;
  wire n5394;
  wire n5396;
  wire n5398;
  wire n5399;
  wire n5401;
  wire n5403;
  wire [1:0] n5404;
  wire [3:0] n5405;
  wire [1:0] n5406;
  wire n5407;
  wire n5408;
  wire n5409;
  wire n5410;
  wire n5411;
  wire n5412;
  wire n5413;
  wire n5414;
  wire n5415;
  wire n5416;
  wire n5417;
  wire n5418;
  wire n5419;
  wire n5420;
  wire n5421;
  wire n5422;
  wire n5423;
  wire [3:0] n5424;
  wire [3:0] n5425;
  wire n5426;
  wire [1:0] n5427;
  wire n5428;
  wire n5429;
  wire [2:0] n5430;
  wire n5432;
  wire n5434;
  wire [2:0] n5436;
  wire [6:0] n5437;
  wire n5439;
  wire [6:0] n5440;
  reg n5441;
  reg [1:0] n5442;
  reg [1:0] n5443;
  reg n5444;
  reg n5445;
  reg n5447;
  reg n5448;
  reg n5450;
  reg n5452;
  reg n5454;
  reg n5456;
  reg n5458;
  reg n5460;
  reg n5462;
  reg n5464;
  reg [5:0] n5465;
  reg n5467;
  reg n5468;
  reg n5470;
  reg n5472;
  reg n5474;
  reg n5476;
  reg n5478;
  reg n5480;
  reg n5482;
  wire n5483;
  reg n5484;
  wire n5485;
  reg n5486;
  wire n5487;
  reg n5488;
  wire n5489;
  reg n5490;
  wire n5491;
  reg n5492;
  wire n5493;
  reg n5494;
  wire n5495;
  reg n5496;
  wire n5497;
  reg n5498;
  wire n5499;
  reg n5500;
  wire n5501;
  reg n5502;
  wire n5503;
  reg n5504;
  wire n5505;
  reg n5506;
  wire n5507;
  wire n5508;
  reg n5509;
  wire n5510;
  wire n5511;
  reg n5512;
  wire n5513;
  reg n5514;
  wire n5515;
  reg n5516;
  wire n5517;
  reg n5518;
  wire n5519;
  reg n5520;
  wire [3:0] n5521;
  reg [3:0] n5522;
  reg [1:0] n5523;
  reg [1:0] n5524;
  wire n5525;
  reg n5526;
  wire n5527;
  reg n5528;
  wire n5529;
  reg n5530;
  reg n5531;
  wire n5532;
  reg n5533;
  reg n5535;
  wire n5536;
  reg n5538;
  wire n5539;
  reg n5541;
  reg n5543;
  reg n5545;
  reg n5547;
  reg n5549;
  reg n5551;
  reg n5553;
  reg n5555;
  reg n5557;
  wire [1:0] n5558;
  reg [1:0] n5560;
  wire n5561;
  reg n5563;
  reg n5565;
  reg [6:0] n5566;
  wire n5567;
  wire [1:0] n5568;
  wire [1:0] n5569;
  wire n5570;
  wire n5571;
  wire n5573;
  wire n5574;
  wire n5576;
  wire n5578;
  wire n5579;
  wire n5580;
  wire n5581;
  wire n5583;
  wire n5585;
  wire n5587;
  wire n5588;
  wire [5:0] n5589;
  wire n5591;
  wire n5592;
  wire n5593;
  wire n5595;
  wire n5597;
  wire n5599;
  wire n5600;
  wire n5602;
  wire n5603;
  wire [3:0] n5604;
  wire [9:0] n5605;
  wire [4:0] n5606;
  wire [1:0] n5607;
  wire n5608;
  wire n5609;
  wire n5610;
  wire n5611;
  wire n5612;
  wire n5613;
  wire n5614;
  wire n5615;
  wire n5616;
  wire n5617;
  wire n5618;
  wire n5619;
  wire n5620;
  wire n5621;
  wire n5622;
  wire n5623;
  wire n5624;
  wire n5625;
  wire [2:0] n5626;
  wire n5627;
  wire [2:0] n5628;
  wire [2:0] n5629;
  wire n5630;
  wire n5631;
  wire [4:0] n5632;
  wire [4:0] n5633;
  wire [4:0] n5634;
  wire n5635;
  wire n5636;
  wire [3:0] n5637;
  wire [3:0] n5638;
  wire [3:0] n5639;
  wire n5640;
  wire [4:0] n5641;
  wire [4:0] n5642;
  wire n5643;
  wire n5644;
  wire n5645;
  wire n5646;
  wire n5647;
  wire [1:0] n5648;
  wire [1:0] n5649;
  wire [1:0] n5650;
  wire [1:0] n5651;
  wire [2:0] n5652;
  wire n5653;
  wire [1:0] n5655;
  wire [1:0] n5657;
  wire n5658;
  wire n5660;
  wire n5662;
  wire n5664;
  wire n5666;
  wire n5668;
  wire n5670;
  wire [1:0] n5671;
  wire [1:0] n5673;
  wire n5674;
  wire n5675;
  wire n5676;
  wire [6:0] n5677;
  wire n5679;
  wire [1:0] n5680;
  wire n5682;
  wire [2:0] n5683;
  wire n5685;
  wire n5689;
  wire n5690;
  wire n5691;
  wire [6:0] n5693;
  wire [2:0] n5694;
  wire n5696;
  wire [1:0] n5697;
  wire n5699;
  wire [2:0] n5700;
  wire n5702;
  wire n5703;
  wire n5704;
  wire n5705;
  wire [1:0] n5706;
  wire n5708;
  wire n5709;
  wire n5711;
  wire n5712;
  wire [6:0] n5714;
  wire [1:0] n5716;
  wire [1:0] n5717;
  wire n5718;
  wire n5719;
  wire n5720;
  wire n5721;
  wire n5724;
  wire n5727;
  wire [1:0] n5728;
  wire n5731;
  wire n5733;
  wire n5735;
  wire n5736;
  wire n5737;
  wire [2:0] n5738;
  wire n5740;
  wire [1:0] n5741;
  wire n5743;
  wire n5744;
  wire n5746;
  wire n5748;
  wire n5749;
  wire n5750;
  wire n5751;
  wire n5753;
  wire [1:0] n5754;
  wire n5756;
  wire n5759;
  wire n5760;
  wire [1:0] n5762;
  wire n5765;
  wire n5768;
  wire n5771;
  wire n5774;
  wire n5776;
  wire n5778;
  wire n5779;
  wire [1:0] n5780;
  wire n5781;
  wire n5783;
  wire n5784;
  wire n5786;
  wire n5787;
  wire n5789;
  wire n5790;
  wire n5792;
  wire n5794;
  wire n5795;
  wire n5796;
  wire [1:0] n5797;
  wire [1:0] n5798;
  wire n5800;
  wire n5802;
  wire n5804;
  wire n5806;
  wire n5808;
  wire n5810;
  wire n5812;
  wire n5813;
  wire n5815;
  wire n5817;
  wire [6:0] n5818;
  wire [4:0] n5819;
  wire n5821;
  wire [2:0] n5822;
  wire n5824;
  wire [1:0] n5825;
  wire n5827;
  wire n5828;
  wire n5829;
  wire [2:0] n5830;
  wire n5832;
  wire n5834;
  wire n5835;
  wire n5836;
  wire n5838;
  wire n5839;
  wire [1:0] n5843;
  wire n5845;
  wire n5848;
  wire n5851;
  wire n5854;
  wire n5857;
  wire n5860;
  wire n5862;
  wire n5864;
  wire [1:0] n5865;
  wire [1:0] n5867;
  wire n5869;
  wire n5871;
  wire n5872;
  wire [1:0] n5873;
  wire [1:0] n5874;
  wire n5876;
  wire n5877;
  wire n5878;
  wire n5880;
  wire n5881;
  wire n5882;
  wire n5883;
  wire n5884;
  wire n5886;
  wire n5887;
  wire n5888;
  wire n5889;
  wire [1:0] n5891;
  wire n5893;
  wire n5895;
  wire n5896;
  wire [6:0] n5897;
  wire n5899;
  wire n5901;
  wire [3:0] n5902;
  wire n5904;
  wire [7:0] n5906;
  wire n5908;
  wire [7:0] n5910;
  wire n5912;
  wire [1:0] n5914;
  wire n5917;
  wire [6:0] n5920;
  wire [1:0] n5921;
  wire n5923;
  wire n5924;
  wire [6:0] n5926;
  wire [7:0] n5927;
  wire n5929;
  wire [7:0] n5931;
  wire n5933;
  wire [1:0] n5935;
  wire [1:0] n5936;
  wire n5937;
  wire [1:0] n5938;
  wire n5940;
  wire n5942;
  wire n5943;
  wire n5944;
  wire n5945;
  wire [6:0] n5947;
  wire [1:0] n5948;
  wire n5949;
  wire n5951;
  wire n5953;
  wire n5954;
  wire [6:0] n5955;
  wire n5957;
  wire n5958;
  wire n5959;
  wire [1:0] n5964;
  wire n5967;
  wire n5970;
  wire n5973;
  wire [1:0] n5974;
  wire [1:0] n5976;
  wire n5978;
  wire n5980;
  wire [1:0] n5981;
  wire n5983;
  wire [2:0] n5984;
  wire n5986;
  wire n5988;
  wire [3:0] n5989;
  wire n5991;
  wire [1:0] n5992;
  wire n5994;
  wire n5995;
  wire n5996;
  wire [1:0] n5997;
  wire n5999;
  wire n6002;
  wire n6004;
  wire n6005;
  wire [1:0] n6006;
  wire n6008;
  wire n6009;
  wire n6010;
  wire [1:0] n6012;
  wire [6:0] n6014;
  wire n6015;
  wire n6016;
  wire n6017;
  wire n6020;
  wire [1:0] n6021;
  wire n6023;
  wire n6024;
  wire n6025;
  wire n6028;
  wire [1:0] n6030;
  wire n6031;
  wire n6033;
  wire n6036;
  wire n6038;
  wire n6041;
  wire n6044;
  wire n6047;
  wire n6049;
  wire n6050;
  wire n6051;
  wire [1:0] n6052;
  wire n6054;
  wire n6055;
  wire [1:0] n6056;
  wire n6058;
  wire [1:0] n6062;
  wire n6064;
  wire [1:0] n6065;
  wire n6067;
  wire n6068;
  wire [1:0] n6071;
  wire n6073;
  wire [1:0] n6078;
  wire n6080;
  wire n6082;
  wire n6083;
  wire n6084;
  wire [1:0] n6085;
  wire n6087;
  wire [1:0] n6090;
  wire n6094;
  wire n6095;
  wire n6096;
  wire n6097;
  wire [6:0] n6099;
  wire n6101;
  wire [6:0] n6103;
  wire [1:0] n6104;
  wire n6107;
  wire n6110;
  wire n6111;
  wire n6113;
  wire n6115;
  wire n6117;
  wire [6:0] n6118;
  wire [1:0] n6119;
  wire n6120;
  wire n6122;
  wire n6125;
  wire n6127;
  wire n6128;
  wire n6131;
  wire n6134;
  wire n6136;
  wire n6137;
  wire n6138;
  wire n6140;
  wire [1:0] n6141;
  wire n6143;
  wire n6145;
  wire [1:0] n6147;
  wire [6:0] n6148;
  wire [1:0] n6149;
  wire [1:0] n6150;
  wire n6152;
  wire n6154;
  wire n6156;
  wire n6157;
  wire n6159;
  wire n6161;
  wire n6164;
  wire n6165;
  wire n6166;
  wire n6167;
  wire n6168;
  wire n6169;
  wire n6170;
  wire n6171;
  wire n6172;
  wire n6174;
  wire n6176;
  wire n6178;
  wire n6180;
  wire [1:0] n6182;
  wire [6:0] n6183;
  wire [1:0] n6184;
  wire n6186;
  wire n6187;
  wire n6188;
  wire [2:0] n6189;
  wire n6191;
  wire n6192;
  wire [3:0] n6193;
  wire n6195;
  wire [1:0] n6196;
  wire n6198;
  wire n6199;
  wire n6200;
  wire n6201;
  wire [1:0] n6202;
  wire n6204;
  wire n6205;
  wire [2:0] n6206;
  wire n6208;
  wire [1:0] n6209;
  wire n6211;
  wire n6212;
  wire n6213;
  wire n6214;
  wire n6215;
  wire n6219;
  wire n6222;
  wire n6225;
  wire n6227;
  wire [1:0] n6228;
  wire [1:0] n6229;
  wire n6231;
  wire n6233;
  wire n6235;
  wire n6236;
  wire n6237;
  wire n6238;
  wire n6240;
  wire n6242;
  wire n6243;
  wire n6244;
  wire n6245;
  wire n6246;
  wire n6248;
  wire n6249;
  wire n6250;
  wire n6252;
  wire n6254;
  wire n6256;
  wire n6258;
  wire n6260;
  wire [1:0] n6262;
  wire [6:0] n6263;
  wire [1:0] n6264;
  wire [1:0] n6265;
  wire n6266;
  wire n6268;
  wire n6270;
  wire n6271;
  wire n6272;
  wire n6273;
  wire n6274;
  wire n6275;
  wire n6277;
  wire n6279;
  wire n6281;
  wire n6282;
  wire n6283;
  wire n6284;
  wire n6285;
  wire n6286;
  wire n6287;
  wire n6288;
  wire n6289;
  wire n6291;
  wire n6293;
  wire n6295;
  wire n6297;
  wire n6298;
  wire [1:0] n6300;
  wire [6:0] n6301;
  wire n6303;
  wire [5:0] n6304;
  wire n6306;
  wire n6307;
  wire n6308;
  wire [1:0] n6309;
  wire n6311;
  wire n6312;
  wire [3:0] n6313;
  wire n6315;
  wire [1:0] n6316;
  wire n6318;
  wire n6319;
  wire n6320;
  wire n6321;
  wire [2:0] n6322;
  wire n6324;
  wire [1:0] n6325;
  wire n6327;
  wire n6328;
  wire n6329;
  wire n6330;
  wire n6331;
  wire n6333;
  wire n6334;
  wire n6336;
  wire n6337;
  wire [1:0] n6338;
  wire n6340;
  wire n6341;
  wire n6342;
  wire [1:0] n6344;
  wire n6346;
  wire n6349;
  wire n6353;
  wire n6356;
  wire n6357;
  wire [1:0] n6358;
  wire n6360;
  wire n6361;
  wire n6364;
  wire n6367;
  wire n6368;
  wire n6370;
  wire n6373;
  wire n6375;
  wire n6377;
  wire n6379;
  wire n6381;
  wire n6382;
  wire n6383;
  wire n6385;
  wire n6386;
  wire n6388;
  wire n6390;
  wire n6392;
  wire n6394;
  wire n6397;
  wire n6400;
  wire n6403;
  wire n6405;
  wire n6407;
  wire n6409;
  wire n6411;
  wire n6413;
  wire n6415;
  wire n6417;
  wire n6419;
  wire n6420;
  wire n6422;
  wire [1:0] n6423;
  wire n6425;
  wire [3:0] n6426;
  wire n6428;
  wire [1:0] n6429;
  wire n6431;
  wire n6432;
  wire n6433;
  wire n6434;
  wire [1:0] n6437;
  wire n6439;
  wire n6441;
  wire n6444;
  wire n6446;
  wire n6449;
  wire n6452;
  wire n6455;
  wire n6457;
  wire n6459;
  wire n6461;
  wire n6463;
  wire n6465;
  wire n6468;
  wire n6471;
  wire n6474;
  wire n6475;
  wire n6476;
  wire n6478;
  wire n6480;
  wire n6481;
  wire [2:0] n6482;
  wire n6484;
  wire [2:0] n6486;
  wire n6488;
  wire n6490;
  wire [1:0] n6494;
  wire n6495;
  wire n6496;
  wire n6497;
  wire n6498;
  wire [6:0] n6500;
  wire [2:0] n6503;
  wire n6505;
  wire [1:0] n6506;
  wire n6508;
  wire n6509;
  wire n6513;
  wire n6516;
  wire n6519;
  wire n6522;
  wire n6524;
  wire n6525;
  wire n6527;
  wire n6529;
  wire n6531;
  wire n6533;
  wire n6534;
  wire n6536;
  wire n6537;
  wire n6538;
  wire n6539;
  wire n6541;
  wire n6543;
  wire n6545;
  wire n6546;
  wire [5:0] n6547;
  wire n6549;
  wire [3:0] n6550;
  wire n6552;
  wire [1:0] n6553;
  wire n6555;
  wire n6556;
  wire n6557;
  wire n6562;
  wire n6565;
  wire n6568;
  wire n6571;
  wire n6572;
  wire n6573;
  wire n6575;
  wire n6576;
  wire n6577;
  wire n6578;
  wire n6579;
  wire n6580;
  wire n6581;
  wire n6583;
  wire n6584;
  wire n6585;
  wire [1:0] n6586;
  wire n6587;
  wire n6589;
  wire n6590;
  wire n6591;
  wire n6593;
  wire n6594;
  wire n6595;
  wire [1:0] n6596;
  wire n6598;
  wire n6600;
  wire n6602;
  wire n6604;
  wire n6605;
  wire n6606;
  wire n6607;
  wire n6609;
  wire n6610;
  wire n6611;
  wire n6612;
  wire n6613;
  wire n6614;
  wire [1:0] n6615;
  wire n6616;
  wire n6618;
  wire n6619;
  wire n6620;
  wire n6622;
  wire n6624;
  wire [6:0] n6625;
  wire n6627;
  wire [1:0] n6628;
  wire n6630;
  wire [2:0] n6631;
  wire n6633;
  wire n6635;
  wire [3:0] n6636;
  wire n6638;
  wire [1:0] n6639;
  wire n6641;
  wire n6642;
  wire n6643;
  wire [1:0] n6644;
  wire n6646;
  wire n6649;
  wire n6651;
  wire n6652;
  wire [1:0] n6653;
  wire n6655;
  wire n6656;
  wire n6657;
  wire n6661;
  wire n6663;
  wire [1:0] n6665;
  wire n6667;
  wire n6668;
  wire n6669;
  wire n6672;
  wire [1:0] n6675;
  wire [1:0] n6677;
  wire n6679;
  wire n6682;
  wire n6684;
  wire n6687;
  wire n6690;
  wire n6693;
  wire n6695;
  wire n6697;
  wire n6699;
  wire n6700;
  wire [1:0] n6701;
  wire n6703;
  wire n6704;
  wire [1:0] n6705;
  wire n6707;
  wire [3:0] n6710;
  wire n6712;
  wire [4:0] n6713;
  wire n6715;
  wire n6716;
  wire n6720;
  wire n6721;
  wire n6722;
  wire n6725;
  wire n6728;
  wire [1:0] n6730;
  wire n6733;
  wire [1:0] n6735;
  wire n6736;
  wire n6738;
  wire n6740;
  wire n6742;
  wire n6745;
  wire n6748;
  wire n6749;
  wire n6750;
  wire n6751;
  wire n6752;
  wire n6753;
  wire n6754;
  wire [1:0] n6755;
  wire [1:0] n6756;
  wire n6758;
  wire n6760;
  wire n6762;
  wire n6764;
  wire n6766;
  wire n6769;
  wire n6770;
  wire n6771;
  wire n6772;
  wire n6773;
  wire n6774;
  wire n6775;
  wire n6777;
  wire n6779;
  wire [1:0] n6780;
  wire n6782;
  wire n6783;
  wire n6784;
  wire [2:0] n6785;
  wire n6787;
  wire n6788;
  wire [3:0] n6789;
  wire n6791;
  wire [1:0] n6792;
  wire n6794;
  wire n6795;
  wire n6796;
  wire n6797;
  wire [1:0] n6798;
  wire n6800;
  wire n6801;
  wire [2:0] n6802;
  wire n6804;
  wire [1:0] n6805;
  wire n6807;
  wire n6808;
  wire n6809;
  wire n6810;
  wire n6811;
  wire n6815;
  wire n6818;
  wire n6821;
  wire n6823;
  wire [1:0] n6824;
  wire [1:0] n6825;
  wire n6827;
  wire n6829;
  wire n6831;
  wire n6832;
  wire n6833;
  wire n6835;
  wire n6837;
  wire n6838;
  wire n6839;
  wire n6840;
  wire n6841;
  wire n6842;
  wire n6843;
  wire n6845;
  wire n6847;
  wire n6849;
  wire [1:0] n6850;
  wire [1:0] n6851;
  wire n6853;
  wire n6855;
  wire n6857;
  wire n6859;
  wire n6860;
  wire n6861;
  wire n6862;
  wire n6864;
  wire n6866;
  wire n6868;
  wire n6869;
  wire n6870;
  wire n6871;
  wire n6872;
  wire n6873;
  wire n6874;
  wire n6876;
  wire n6878;
  wire n6880;
  wire n6882;
  wire n6884;
  wire n6886;
  wire n6888;
  wire [1:0] n6889;
  wire n6891;
  wire n6892;
  wire n6893;
  wire [1:0] n6894;
  wire n6896;
  wire [2:0] n6897;
  wire n6899;
  wire [1:0] n6900;
  wire n6902;
  wire n6903;
  wire n6904;
  wire [1:0] n6906;
  wire [1:0] n6909;
  wire n6912;
  wire [1:0] n6913;
  wire n6916;
  wire n6919;
  wire n6922;
  wire n6924;
  wire n6926;
  wire n6927;
  wire n6928;
  wire n6930;
  wire n6932;
  wire [1:0] n6933;
  wire n6935;
  wire [2:0] n6936;
  wire n6938;
  wire n6939;
  wire [2:0] n6940;
  wire n6942;
  wire n6943;
  wire [2:0] n6944;
  wire n6946;
  wire [2:0] n6947;
  wire n6949;
  wire n6950;
  wire [2:0] n6951;
  wire n6953;
  wire n6954;
  wire [2:0] n6955;
  wire n6957;
  wire [1:0] n6958;
  wire n6960;
  wire n6961;
  wire n6962;
  wire n6963;
  wire n6964;
  wire [1:0] n6965;
  wire n6967;
  wire [2:0] n6968;
  wire n6970;
  wire n6971;
  wire [2:0] n6972;
  wire n6974;
  wire n6975;
  wire [2:0] n6976;
  wire n6978;
  wire [2:0] n6979;
  wire n6981;
  wire n6982;
  wire [2:0] n6983;
  wire n6985;
  wire n6986;
  wire [3:0] n6987;
  wire n6989;
  wire n6990;
  wire n6991;
  wire n6992;
  wire n6995;
  wire n6996;
  wire n6997;
  wire n6998;
  wire [6:0] n7000;
  wire n7002;
  wire n7003;
  wire n7004;
  wire n7005;
  wire n7008;
  wire [2:0] n7009;
  wire n7011;
  wire n7014;
  wire [2:0] n7015;
  wire n7017;
  wire [2:0] n7018;
  wire n7020;
  wire n7021;
  wire [2:0] n7022;
  wire n7024;
  wire n7025;
  wire [2:0] n7026;
  wire n7028;
  wire n7029;
  wire n7032;
  wire [2:0] n7033;
  wire n7035;
  wire [2:0] n7036;
  wire n7038;
  wire n7039;
  wire [2:0] n7040;
  wire n7042;
  wire n7043;
  wire n7046;
  wire [1:0] n7047;
  wire n7049;
  wire [2:0] n7050;
  wire n7052;
  wire n7054;
  wire n7055;
  wire [1:0] n7058;
  wire n7061;
  wire n7064;
  wire n7065;
  wire n7066;
  wire n7067;
  wire n7069;
  wire n7071;
  wire n7073;
  wire n7074;
  wire n7075;
  wire [1:0] n7077;
  wire n7078;
  wire [1:0] n7082;
  wire n7084;
  wire n7086;
  wire n7087;
  wire n7088;
  wire n7089;
  wire [6:0] n7091;
  wire [2:0] n7092;
  wire n7094;
  wire n7097;
  wire n7100;
  wire [2:0] n7101;
  wire n7103;
  wire [2:0] n7104;
  wire n7106;
  wire n7107;
  wire [2:0] n7108;
  wire n7110;
  wire n7111;
  wire n7113;
  wire n7115;
  wire n7117;
  wire n7118;
  wire [1:0] n7119;
  wire n7121;
  wire n7124;
  wire n7126;
  wire n7128;
  wire n7130;
  wire n7132;
  wire n7135;
  wire n7138;
  wire n7139;
  wire n7140;
  wire n7141;
  wire n7142;
  wire n7143;
  wire n7144;
  wire n7145;
  wire n7146;
  wire [1:0] n7147;
  wire n7149;
  wire n7151;
  wire [1:0] n7153;
  wire [6:0] n7154;
  wire n7155;
  wire [1:0] n7156;
  wire n7157;
  wire n7159;
  wire n7161;
  wire n7163;
  wire n7165;
  wire n7167;
  wire n7168;
  wire n7169;
  wire n7170;
  wire n7172;
  wire n7173;
  wire n7174;
  wire n7175;
  wire n7176;
  wire n7177;
  wire n7178;
  wire n7179;
  wire n7180;
  wire n7181;
  wire n7183;
  wire [1:0] n7185;
  wire n7187;
  wire [6:0] n7188;
  wire n7189;
  wire n7190;
  wire n7192;
  wire n7194;
  wire [1:0] n7196;
  wire n7198;
  wire [2:0] n7200;
  wire [2:0] n7201;
  wire n7203;
  wire n7206;
  wire [1:0] n7208;
  wire [3:0] n7209;
  wire [3:0] n7210;
  wire [3:0] n7211;
  wire n7212;
  wire n7213;
  wire [6:0] n7215;
  wire n7216;
  wire [3:0] n7217;
  wire [3:0] n7218;
  wire n7220;
  wire n7221;
  wire [1:0] n7223;
  wire n7225;
  wire [1:0] n7226;
  wire n7228;
  wire n7230;
  wire n7232;
  wire n7233;
  wire n7235;
  wire n7236;
  wire n7237;
  wire [1:0] n7238;
  wire n7241;
  wire n7243;
  wire n7245;
  wire n7247;
  wire n7249;
  wire n7251;
  wire n7253;
  wire [1:0] n7254;
  wire [3:0] n7255;
  wire [3:0] n7256;
  wire n7258;
  wire n7260;
  wire n7262;
  wire n7263;
  wire n7264;
  wire n7265;
  wire n7266;
  wire n7267;
  wire n7268;
  wire n7269;
  wire n7270;
  wire n7271;
  wire n7272;
  wire n7274;
  wire n7276;
  wire n7277;
  wire [1:0] n7279;
  wire n7280;
  wire [6:0] n7281;
  wire n7283;
  wire n7284;
  wire [2:0] n7285;
  wire n7287;
  wire n7288;
  wire [1:0] n7289;
  wire n7291;
  wire [2:0] n7292;
  wire n7294;
  wire n7295;
  wire [2:0] n7296;
  wire n7298;
  wire [1:0] n7299;
  wire n7301;
  wire n7302;
  wire n7303;
  wire [2:0] n7304;
  wire n7306;
  wire n7307;
  wire n7308;
  wire [1:0] n7309;
  wire n7311;
  wire n7312;
  wire n7315;
  wire n7318;
  wire n7320;
  wire n7323;
  wire n7325;
  wire n7328;
  wire n7331;
  wire n7333;
  wire n7334;
  wire n7335;
  wire n7337;
  wire n7339;
  wire n7341;
  wire n7342;
  wire [2:0] n7343;
  wire n7345;
  wire n7346;
  wire [1:0] n7347;
  wire n7349;
  wire [2:0] n7350;
  wire n7352;
  wire n7353;
  wire [2:0] n7354;
  wire n7356;
  wire [1:0] n7357;
  wire n7359;
  wire [2:0] n7360;
  wire n7362;
  wire n7363;
  wire n7364;
  wire n7365;
  wire [4:0] n7366;
  wire n7368;
  wire [2:0] n7369;
  wire n7371;
  wire [2:0] n7372;
  wire n7374;
  wire n7375;
  wire [2:0] n7376;
  wire n7378;
  wire n7381;
  wire n7384;
  wire n7386;
  wire n7389;
  wire n7391;
  wire n7394;
  wire n7397;
  wire n7399;
  wire n7400;
  wire n7401;
  wire n7403;
  wire n7405;
  wire n7407;
  wire n7409;
  wire n7411;
  wire n7413;
  wire n7415;
  wire n7417;
  wire n7419;
  wire n7420;
  wire n7421;
  wire n7422;
  wire n7424;
  wire [12:0] n7425;
  reg n7426;
  reg [1:0] n7428;
  reg [1:0] n7429;
  reg [1:0] n7430;
  reg n7431;
  reg n7433;
  reg n7435;
  reg n7437;
  reg n7440;
  reg n7442;
  reg n7444;
  reg n7447;
  reg n7450;
  reg n7453;
  reg n7456;
  reg n7459;
  reg n7462;
  reg n7465;
  reg n7468;
  reg n7471;
  reg [1:0] n7473;
  wire [3:0] n7474;
  wire [3:0] n7475;
  reg [3:0] n7476;
  wire [1:0] n7477;
  wire [1:0] n7478;
  reg [1:0] n7479;
  reg n7482;
  reg n7484;
  reg n7487;
  reg n7490;
  reg n7494;
  reg n7497;
  reg n7500;
  reg n7503;
  reg n7509;
  reg n7512;
  reg n7515;
  reg n7518;
  reg n7521;
  reg n7524;
  wire n7526;
  reg n7527;
  wire [2:0] n7528;
  reg [2:0] n7529;
  wire n7530;
  reg n7531;
  wire n7532;
  reg n7533;
  wire n7534;
  reg n7535;
  wire n7536;
  reg n7537;
  wire n7538;
  reg n7539;
  wire n7540;
  reg n7541;
  wire n7542;
  reg n7543;
  reg n7544;
  wire n7545;
  reg n7546;
  wire n7547;
  reg n7548;
  wire n7549;
  wire n7550;
  reg n7551;
  wire n7552;
  wire n7553;
  reg n7554;
  wire n7555;
  reg n7556;
  wire n7557;
  wire n7558;
  wire n7559;
  reg n7560;
  wire n7561;
  wire n7562;
  wire n7563;
  reg n7564;
  wire n7565;
  wire n7566;
  reg n7567;
  wire n7568;
  wire n7569;
  reg n7570;
  wire n7571;
  reg n7572;
  wire [1:0] n7573;
  wire [1:0] n7574;
  reg [1:0] n7575;
  wire n7576;
  wire n7577;
  reg n7578;
  wire n7579;
  wire n7580;
  reg n7581;
  wire n7582;
  wire n7583;
  wire n7584;
  reg n7585;
  wire n7586;
  wire n7587;
  reg n7588;
  wire [3:0] n7589;
  reg [3:0] n7590;
  wire n7591;
  reg n7592;
  wire n7593;
  wire [4:0] n7594;
  reg [4:0] n7595;
  wire n7596;
  reg n7597;
  wire n7598;
  reg n7599;
  wire n7600;
  reg n7601;
  wire n7602;
  wire n7603;
  reg n7604;
  wire n7605;
  reg n7606;
  wire n7607;
  reg n7608;
  wire n7609;
  reg n7610;
  wire n7611;
  reg n7612;
  wire n7613;
  reg n7614;
  wire [15:0] n7617;
  wire n7618;
  wire n7619;
  wire [3:0] n7624;
  wire n7626;
  wire n7630;
  wire n7641;
  wire n7642;
  wire n7643;
  wire n7647;
  wire n7651;
  reg n7653;
  wire n7654;
  reg n7656;
  wire n7657;
  reg n7659;
  wire n7660;
  wire n7661;
  reg n7663;
  wire n7664;
  reg n7666;
  wire n7667;
  reg n7669;
  wire n7670;
  wire n7671;
  reg n7673;
  wire n7674;
  wire n7675;
  reg n7677;
  wire n7678;
  reg n7680;
  reg n7682;
  reg n7684;
  reg n7686;
  reg n7688;
  reg n7690;
  reg n7692;
  reg n7694;
  reg n7696;
  reg n7698;
  reg n7700;
  reg n7702;
  reg n7704;
  reg n7706;
  reg [1:0] n7708;
  reg n7710;
  reg n7712;
  reg [1:0] n7714;
  reg [1:0] n7716;
  reg n7718;
  reg n7720;
  localparam [88:0] n7721 = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [2:0] n7740;
  wire n7744;
  wire n7746;
  wire [31:0] n7751;
  wire [6:0] n7753;
  wire [1:0] n7756;
  wire [5:0] n7757;
  reg [6:0] n7758;
  wire n7759;
  wire n7760;
  wire n7761;
  wire n7762;
  wire [1:0] n7763;
  wire n7765;
  wire n7766;
  wire n7767;
  wire n7769;
  wire n7770;
  wire n7772;
  wire n7774;
  wire n7776;
  wire n7778;
  wire n7779;
  wire n7781;
  wire n7782;
  wire n7783;
  wire n7784;
  wire n7785;
  wire n7786;
  wire n7787;
  wire n7789;
  wire n7790;
  wire n7791;
  wire n7794;
  wire [2:0] n7795;
  wire n7797;
  wire n7799;
  wire [1:0] n7803;
  wire n7805;
  wire n7806;
  wire n7807;
  wire n7808;
  wire [6:0] n7810;
  wire n7812;
  wire n7813;
  wire n7815;
  wire n7816;
  wire n7817;
  wire n7818;
  wire n7819;
  wire n7820;
  wire n7821;
  wire n7823;
  wire n7825;
  wire n7826;
  wire n7827;
  wire n7828;
  wire n7829;
  wire n7830;
  wire n7831;
  wire n7832;
  wire n7833;
  wire n7834;
  wire n7835;
  wire n7837;
  wire n7838;
  wire n7840;
  wire n7842;
  wire [6:0] n7843;
  wire n7844;
  wire [6:0] n7846;
  wire n7852;
  wire n7855;
  wire n7858;
  wire n7859;
  wire n7860;
  wire n7862;
  wire n7863;
  wire n7864;
  wire n7866;
  wire n7867;
  wire n7869;
  wire n7870;
  wire n7872;
  wire n7874;
  wire n7875;
  wire n7876;
  wire n7877;
  wire n7878;
  wire n7880;
  wire [1:0] n7882;
  wire n7883;
  wire [1:0] n7885;
  wire n7888;
  wire n7891;
  wire n7892;
  wire n7893;
  wire n7894;
  wire n7895;
  wire [6:0] n7898;
  wire n7900;
  wire n7903;
  wire n7904;
  wire n7907;
  wire n7908;
  wire n7909;
  wire n7910;
  wire n7911;
  wire n7912;
  wire [1:0] n7914;
  wire n7916;
  wire [6:0] n7919;
  wire [1:0] n7920;
  wire n7922;
  wire [1:0] n7926;
  wire n7929;
  wire n7931;
  wire n7932;
  wire n7933;
  wire [6:0] n7935;
  wire [1:0] n7937;
  wire n7939;
  wire n7940;
  wire n7941;
  wire n7942;
  wire n7943;
  wire [6:0] n7944;
  wire n7946;
  wire n7949;
  wire n7951;
  wire n7952;
  wire n7953;
  wire n7955;
  wire [1:0] n7957;
  wire n7958;
  wire n7960;
  wire n7961;
  wire n7964;
  wire n7965;
  wire n7966;
  wire n7967;
  wire n7968;
  wire [1:0] n7972;
  wire n7974;
  wire n7975;
  wire n7976;
  wire [6:0] n7978;
  wire n7980;
  wire n7982;
  wire n7983;
  wire n7984;
  wire n7986;
  wire n7987;
  wire n7988;
  wire n7990;
  wire n7991;
  wire n7993;
  wire n7995;
  wire n7996;
  wire n7997;
  wire n7998;
  wire n8000;
  wire [1:0] n8002;
  wire n8003;
  wire [1:0] n8005;
  wire n8008;
  wire n8011;
  wire n8012;
  wire n8013;
  wire n8014;
  wire [6:0] n8017;
  wire n8019;
  wire n8022;
  wire n8023;
  wire n8026;
  wire n8027;
  wire n8028;
  wire n8029;
  wire n8030;
  wire n8031;
  wire [1:0] n8033;
  wire n8035;
  wire [6:0] n8038;
  wire [1:0] n8039;
  wire n8041;
  wire [1:0] n8046;
  wire n8047;
  wire n8048;
  wire n8049;
  wire [6:0] n8052;
  wire [1:0] n8054;
  wire n8055;
  wire n8056;
  wire n8057;
  wire n8058;
  wire [6:0] n8059;
  wire n8061;
  wire n8065;
  wire n8068;
  wire n8069;
  wire n8070;
  wire n8072;
  wire [1:0] n8074;
  wire n8075;
  wire n8077;
  wire n8079;
  wire n8082;
  wire n8083;
  wire n8084;
  wire n8085;
  wire n8086;
  wire [1:0] n8090;
  wire n8091;
  wire [6:0] n8094;
  wire n8096;
  wire n8098;
  wire n8101;
  wire [6:0] n8103;
  wire n8105;
  wire n8107;
  wire n8108;
  wire n8111;
  wire n8114;
  wire n8116;
  wire n8117;
  wire n8118;
  wire n8120;
  wire n8123;
  wire [6:0] n8125;
  wire n8126;
  wire n8129;
  wire n8131;
  wire n8132;
  wire n8134;
  wire n8140;
  wire n8141;
  wire [1:0] n8142;
  wire n8144;
  wire n8146;
  wire n8147;
  wire [1:0] n8149;
  wire n8152;
  wire n8154;
  wire n8159;
  wire n8161;
  wire [1:0] n8163;
  wire n8166;
  wire n8170;
  wire n8171;
  wire [1:0] n8173;
  wire [6:0] n8175;
  wire n8177;
  wire n8179;
  wire n8180;
  wire n8182;
  wire n8184;
  wire n8186;
  wire n8187;
  wire [1:0] n8194;
  wire n8197;
  wire n8198;
  wire n8199;
  wire n8200;
  wire n8201;
  wire n8202;
  wire n8203;
  wire [6:0] n8205;
  wire n8207;
  wire n8208;
  wire n8211;
  wire n8217;
  wire n8220;
  wire n8221;
  wire n8223;
  wire n8229;
  wire n8232;
  wire n8233;
  wire n8235;
  wire [1:0] n8243;
  wire n8246;
  wire n8248;
  wire n8251;
  wire n8253;
  wire n8254;
  wire n8255;
  wire n8256;
  wire n8257;
  wire n8258;
  wire n8259;
  wire n8260;
  wire n8261;
  wire n8262;
  wire [6:0] n8265;
  wire n8267;
  wire n8271;
  wire n8275;
  wire [15:0] n8276;
  wire n8278;
  wire [2:0] n8279;
  wire n8281;
  wire n8283;
  wire n8285;
  wire n8286;
  wire n8287;
  wire [1:0] n8289;
  wire n8290;
  wire n8291;
  wire [6:0] n8293;
  wire n8295;
  wire n8296;
  wire n8299;
  wire n8300;
  wire [1:0] n8304;
  wire n8305;
  wire [1:0] n8307;
  wire n8308;
  wire n8309;
  wire n8310;
  wire [6:0] n8312;
  wire n8314;
  wire [1:0] n8315;
  wire n8317;
  wire n8319;
  wire n8321;
  wire [2:0] n8322;
  wire n8324;
  wire n8326;
  wire n8331;
  wire [2:0] n8332;
  wire n8334;
  wire n8336;
  wire [1:0] n8338;
  wire n8340;
  wire [1:0] n8343;
  wire n8346;
  wire n8348;
  wire [2:0] n8349;
  wire n8351;
  wire n8353;
  wire n8356;
  wire [2:0] n8357;
  wire n8359;
  wire n8361;
  wire n8364;
  wire n8368;
  wire n8371;
  wire n8374;
  wire n8377;
  wire n8380;
  wire n8383;
  wire n8384;
  wire n8386;
  wire [1:0] n8389;
  wire n8390;
  wire n8391;
  wire [6:0] n8394;
  wire n8396;
  wire n8397;
  wire n8399;
  wire n8402;
  wire [6:0] n8406;
  wire n8408;
  wire n8412;
  wire n8415;
  wire n8418;
  wire n8421;
  wire n8424;
  wire n8425;
  wire n8426;
  wire n8429;
  wire n8430;
  wire n8431;
  wire n8433;
  wire n8435;
  wire n8436;
  wire n8437;
  wire [1:0] n8440;
  wire n8442;
  wire n8443;
  wire [6:0] n8446;
  wire n8448;
  wire n8450;
  wire [3:0] n8451;
  wire n8453;
  wire [1:0] n8457;
  wire [1:0] n8459;
  wire n8461;
  wire n8462;
  wire [6:0] n8465;
  wire n8467;
  wire n8469;
  wire n8471;
  wire n8474;
  wire [11:0] n8476;
  wire n8478;
  wire [11:0] n8479;
  wire n8481;
  wire n8482;
  wire [11:0] n8483;
  wire n8485;
  wire n8486;
  wire [11:0] n8487;
  wire n8489;
  wire n8490;
  wire n8491;
  wire [11:0] n8492;
  wire n8494;
  wire [11:0] n8495;
  wire n8497;
  wire n8498;
  wire [11:0] n8499;
  wire n8501;
  wire n8502;
  wire [11:0] n8503;
  wire n8505;
  wire n8506;
  wire n8507;
  wire n8508;
  wire n8509;
  wire n8510;
  wire n8512;
  wire n8514;
  wire n8516;
  wire n8517;
  wire n8519;
  wire n8523;
  wire n8525;
  wire n8526;
  wire n8527;
  wire [1:0] n8530;
  wire n8532;
  wire n8533;
  wire n8536;
  wire n8537;
  wire n8538;
  wire n8539;
  wire [1:0] n8542;
  wire n8544;
  wire n8545;
  wire n8549;
  wire n8550;
  wire [1:0] n8553;
  wire [1:0] n8555;
  wire [1:0] n8556;
  wire n8557;
  wire n8558;
  wire n8559;
  wire [6:0] n8561;
  wire n8563;
  wire n8564;
  wire n8565;
  wire [1:0] n8568;
  wire n8570;
  wire n8572;
  wire n8573;
  wire n8575;
  wire [5:0] n8578;
  wire n8580;
  wire n8583;
  wire [6:0] n8586;
  wire n8588;
  wire n8589;
  wire n8590;
  wire n8592;
  wire n8594;
  wire n8595;
  wire n8597;
  wire n8599;
  wire [1:0] n8601;
  wire [6:0] n8603;
  wire n8605;
  wire n8607;
  wire n8608;
  wire n8609;
  wire n8610;
  wire n8611;
  wire n8613;
  wire n8618;
  wire n8620;
  wire [15:0] n8621;
  wire n8623;
  wire n8624;
  wire n8625;
  wire n8627;
  wire [15:0] n8628;
  wire n8630;
  wire n8631;
  wire n8634;
  wire [6:0] n8636;
  wire n8639;
  wire n8640;
  wire n8642;
  wire [5:0] n8645;
  wire n8647;
  wire n8650;
  wire [6:0] n8653;
  wire n8655;
  wire n8656;
  wire n8657;
  wire n8658;
  wire n8660;
  wire n8661;
  wire n8662;
  wire n8664;
  wire [1:0] n8667;
  wire n8670;
  wire n8671;
  wire [6:0] n8673;
  wire n8676;
  wire n8677;
  wire n8680;
  wire n8681;
  wire n8684;
  wire [5:0] n8685;
  wire n8687;
  wire [5:0] n8688;
  wire [5:0] n8690;
  wire [5:0] n8691;
  wire n8692;
  wire n8693;
  wire n8695;
  wire n8697;
  wire [80:0] n8698;
  reg n8701;
  reg [1:0] n8714;
  reg [1:0] n8715;
  reg [1:0] n8753;
  reg n8756;
  reg n8759;
  reg n8764;
  reg n8766;
  reg n8776;
  reg n8780;
  reg n8794;
  reg n8796;
  reg n8799;
  reg n8802;
  reg n8805;
  reg n8809;
  reg n8813;
  reg n8816;
  reg n8821;
  reg n8823;
  reg n8828;
  reg n8831;
  reg n8837;
  reg n8841;
  reg n8846;
  wire [5:0] n8847;
  reg [5:0] n8848;
  reg n8852;
  reg n8855;
  reg n8862;
  reg n8864;
  reg n8865;
  reg n8868;
  reg n8870;
  reg n8872;
  reg n8873;
  reg n8874;
  reg n8875;
  reg n8876;
  reg n8877;
  reg n8878;
  wire n8879;
  reg n8880;
  reg n8881;
  reg n8882;
  reg n8883;
  reg n8884;
  reg n8885;
  reg n8886;
  reg n8887;
  reg n8888;
  reg n8889;
  reg n8890;
  reg n8891;
  reg n8892;
  reg n8893;
  wire n8894;
  reg n8895;
  wire n8896;
  reg n8897;
  reg n8898;
  wire n8899;
  reg n8900;
  wire n8901;
  reg n8902;
  reg n8903;
  reg n8904;
  reg n8905;
  reg n8906;
  reg n8907;
  wire n8908;
  reg n8909;
  reg n8910;
  reg n8911;
  reg n8912;
  reg n8913;
  reg n8914;
  wire n8915;
  reg n8916;
  wire n8917;
  reg n8918;
  wire n8919;
  wire [1:0] n8921;
  wire n8923;
  wire [1:0] n8924;
  wire [3:0] n8925;
  wire n8927;
  reg n8928;
  wire [1:0] n8929;
  wire [1:0] n8930;
  reg [6:0] n8971;
  wire n8977;
  wire n8978;
  wire [11:0] n8979;
  wire [2:0] n8980;
  wire n8982;
  wire [2:0] n8983;
  wire n8985;
  wire [3:0] n8986;
  wire n8988;
  wire n8990;
  wire n8992;
  wire n8994;
  wire n8996;
  wire n8998;
  wire [7:0] n8999;
  reg [31:0] n9000;
  reg [3:0] n9001;
  reg [2:0] n9002;
  reg [2:0] n9003;
  wire [31:0] n9004;
  wire [3:0] n9005;
  wire [2:0] n9006;
  wire [2:0] n9007;
  wire [31:0] n9009;
  wire [3:0] n9011;
  wire [2:0] n9012;
  wire [2:0] n9013;
  wire [11:0] n9018;
  wire [31:0] n9020;
  wire n9022;
  wire [31:0] n9024;
  wire n9026;
  wire [3:0] n9028;
  wire [31:0] n9030;
  wire n9032;
  wire n9034;
  wire [3:0] n9035;
  reg [31:0] n9037;
  wire [3:0] n9042;
  wire n9044;
  wire n9046;
  wire n9047;
  wire n9048;
  wire n9049;
  wire n9050;
  wire n9051;
  wire n9053;
  wire n9054;
  wire n9055;
  wire n9056;
  wire n9058;
  wire n9059;
  wire n9060;
  wire n9062;
  wire n9063;
  wire n9065;
  wire n9066;
  wire n9067;
  wire n9069;
  wire n9070;
  wire n9072;
  wire n9073;
  wire n9074;
  wire n9076;
  wire n9077;
  wire n9079;
  wire n9080;
  wire n9081;
  wire n9083;
  wire n9084;
  wire n9086;
  wire n9087;
  wire n9088;
  wire n9089;
  wire n9090;
  wire n9091;
  wire n9092;
  wire n9093;
  wire n9094;
  wire n9095;
  wire n9097;
  wire n9098;
  wire n9099;
  wire n9100;
  wire n9101;
  wire n9102;
  wire n9103;
  wire n9104;
  wire n9105;
  wire n9106;
  wire n9108;
  wire n9109;
  wire n9110;
  wire n9111;
  wire n9112;
  wire n9113;
  wire n9114;
  wire n9115;
  wire n9116;
  wire n9117;
  wire n9118;
  wire n9119;
  wire n9120;
  wire n9121;
  wire n9122;
  wire n9123;
  wire n9125;
  wire n9126;
  wire n9127;
  wire n9128;
  wire n9129;
  wire n9130;
  wire n9131;
  wire n9132;
  wire n9133;
  wire n9134;
  wire n9135;
  wire n9136;
  wire n9138;
  wire [15:0] n9139;
  reg n9142;
  wire n9147;
  wire [15:0] n9148;
  wire n9149;
  wire n9150;
  wire n9151;
  wire n9154;
  wire n9157;
  wire n9160;
  wire n9163;
  wire n9166;
  wire n9169;
  wire n9172;
  wire n9175;
  wire n9178;
  wire n9181;
  wire n9184;
  wire n9187;
  wire n9190;
  wire n9193;
  wire n9196;
  wire n9199;
  wire [15:0] n9200;
  wire n9201;
  reg n9202;
  wire n9203;
  reg n9204;
  wire n9205;
  reg n9206;
  wire n9207;
  reg n9208;
  wire n9209;
  reg n9210;
  wire n9211;
  reg n9212;
  wire n9213;
  reg n9214;
  wire n9215;
  reg n9216;
  wire n9217;
  reg n9218;
  wire n9219;
  reg n9220;
  wire n9221;
  reg n9222;
  wire n9223;
  reg n9224;
  wire n9225;
  reg n9226;
  wire n9227;
  reg n9228;
  wire n9229;
  reg n9230;
  wire n9231;
  reg n9232;
  wire [15:0] n9233;
  wire [15:0] n9234;
  wire [15:0] n9235;
  wire [3:0] n9243;
  wire n9245;
  wire [3:0] n9246;
  wire n9248;
  wire [3:0] n9250;
  wire n9252;
  wire [3:0] n9253;
  wire n9255;
  wire n9258;
  wire [3:0] n9260;
  wire [3:0] n9261;
  wire n9263;
  wire [3:0] n9264;
  wire n9266;
  wire [3:0] n9267;
  wire [1:0] n9269;
  wire n9270;
  wire n9271;
  wire n9272;
  wire n9274;
  wire [3:0] n9275;
  wire n9277;
  wire [3:0] n9278;
  wire [1:0] n9279;
  wire [1:0] n9281;
  localparam [3:0] n9282 = 4'b0000;
  wire [3:0] n9284;
  wire n9286;
  wire [1:0] n9288;
  wire n9290;
  wire n9292;
  wire n9293;
  wire n9295;
  wire n9296;
  wire n9297;
  wire n9298;
  wire n9300;
  wire n9301;
  wire [1:0] n9302;
  wire n9303;
  wire n9304;
  wire n9305;
  wire n9306;
  wire n9307;
  reg n9310;
  wire [3:0] n9311;
  reg [3:0] n9312;
  wire n9313;
  reg n9314;
  reg [31:0] n9315;
  wire [31:0] n9316;
  reg [31:0] n9317;
  wire [31:0] n9318;
  reg [31:0] n9319;
  reg [1:0] n9320;
  reg [1:0] n9321;
  reg n9322;
  reg [15:0] n9323;
  reg [15:0] n9324;
  wire [15:0] n9325;
  reg [15:0] n9326;
  reg [31:0] n9327;
  reg [31:0] n9328;
  reg [15:0] n9329;
  wire [3:0] n9331;
  reg [3:0] n9332;
  wire [31:0] n9333;
  wire [3:0] n9336;
  reg [3:0] n9337;
  wire [3:0] n9338;
  reg [3:0] n9339;
  wire n9340;
  reg n9341;
  wire [31:0] n9342;
  reg [31:0] n9343;
  wire [31:0] n9344;
  reg [31:0] n9345;
  wire n9346;
  reg n9347;
  reg [31:0] n9348;
  wire [31:0] n9349;
  reg [31:0] n9351;
  reg n9352;
  wire [31:0] n9354;
  reg n9355;
  reg [15:0] n9356;
  reg n9357;
  reg n9358;
  reg n9359;
  reg n9360;
  reg n9361;
  reg n9362;
  reg n9363;
  reg [7:0] n9364;
  reg n9365;
  wire n9366;
  reg n9367;
  reg [1:0] n9368;
  reg [5:0] n9369;
  wire n9370;
  reg n9371;
  wire [3:0] n9372;
  reg n9374;
  reg n9375;
  reg n9376;
  reg n9377;
  reg n9378;
  reg n9379;
  reg [7:0] n9380;
  reg n9381;
  reg n9382;
  reg n9383;
  reg n9384;
  wire [31:0] n9385;
  reg [31:0] n9386;
  wire [31:0] n9387;
  reg [31:0] n9388;
  reg [2:0] n9389;
  reg [7:0] n9390;
  reg n9391;
  reg n9392;
  reg n9393;
  reg n9394;
  reg n9395;
  wire [31:0] n9396;
  wire [7:0] n9397;
  reg [7:0] n9398;
  reg [5:0] n9399;
  reg [3:0] n9400;
  reg [5:0] n9401;
  reg n9402;
  reg n9403;
  reg [31:0] n9404;
  reg [31:0] n9405;
  wire [5:0] n9406;
  wire [5:0] n9407;
  reg [5:0] n9408;
  reg [5:0] n9409;
  wire [5:0] n9410;
  reg [31:0] n9411;
  reg [5:0] n9412;
  reg [31:0] n9413;
  reg [3:0] n9414;
  reg [2:0] n9415;
  reg [2:0] n9416;
  wire [88:0] n9417;
  wire [88:0] n9418;
  wire [88:0] n9419;
  reg [88:0] n9420;
  reg [6:0] n9421;
  wire [15:0] n9422;
  reg n9423;
  reg [1:0] n9424;
  wire [2:0] n9425;
  wire [31:0] n9428; // mem_rd
  wire [31:0] n9429; // mem_rd
  assign addr_out = n995; //(module output)
  assign data_write = n9422; //(module output)
  assign nWr = n59; //(module output)
  assign nUDS = n70; //(module output)
  assign nLDS = n71; //(module output)
  assign busstate = state; //(module output)
  assign longword = n37; //(module output)
  assign nResetOut = n63; //(module output)
  assign FC = n9425; //(module output)
  assign clr_berr = n79; //(module output)
  assign skipFetch = n8701; //(module output)
  assign regin_out = regin; //(module output)
  assign CACR_out = cacr; //(module output)
  assign VBR_out = vbr; //(module output)
  /* TG68KdotC_Kernel.vhd:148:16  */
  assign use_vbr_stackframe = n9310; // (signal)
  /* TG68KdotC_Kernel.vhd:150:16  */
  assign syncreset = n9312; // (signal)
  /* TG68KdotC_Kernel.vhd:151:16  */
  assign reset = n9314; // (signal)
  /* TG68KdotC_Kernel.vhd:152:16  */
  assign clkena_lw = n75; // (signal)
  /* TG68KdotC_Kernel.vhd:153:16  */
  assign tg68_pc = n9315; // (signal)
  /* TG68KdotC_Kernel.vhd:154:16  */
  assign tmp_tg68_pc = n9317; // (signal)
  /* TG68KdotC_Kernel.vhd:155:16  */
  assign tg68_pc_add = n1086; // (signal)
  /* TG68KdotC_Kernel.vhd:156:16  */
  assign pc_dataa = n1002; // (signal)
  /* TG68KdotC_Kernel.vhd:157:16  */
  assign pc_datab = n1085; // (signal)
  /* TG68KdotC_Kernel.vhd:158:16  */
  assign memaddr = n9319; // (signal)
  /* TG68KdotC_Kernel.vhd:159:16  */
  assign state = n9320; // (signal)
  /* TG68KdotC_Kernel.vhd:160:16  */
  assign datatype = n8714; // (signal)
  /* TG68KdotC_Kernel.vhd:161:16  */
  assign set_datatype = n8715; // (signal)
  /* TG68KdotC_Kernel.vhd:162:16  */
  assign exe_datatype = n9321; // (signal)
  /* TG68KdotC_Kernel.vhd:163:16  */
  assign setstate = n8753; // (signal)
  /* TG68KdotC_Kernel.vhd:164:16  */
  assign setaddrvalue = n8756; // (signal)
  /* TG68KdotC_Kernel.vhd:165:16  */
  assign addrvalue = n9322; // (signal)
  /* TG68KdotC_Kernel.vhd:167:16  */
  assign opcode = n9323; // (signal)
  /* TG68KdotC_Kernel.vhd:168:16  */
  assign exe_opcode = n9324; // (signal)
  /* TG68KdotC_Kernel.vhd:169:16  */
  assign sndopc = n9326; // (signal)
  /* TG68KdotC_Kernel.vhd:171:16  */
  assign exe_pc = n9327; // (signal)
  /* TG68KdotC_Kernel.vhd:172:16  */
  assign last_opc_pc = n9328; // (signal)
  /* TG68KdotC_Kernel.vhd:173:16  */
  assign last_opc_read = n9329; // (signal)
  /* TG68KdotC_Kernel.vhd:175:16  */
  assign reg_qa = n9429; // (signal)
  /* TG68KdotC_Kernel.vhd:176:16  */
  assign reg_qb = n9428; // (signal)
  /* TG68KdotC_Kernel.vhd:177:16  */
  assign wwrena = n345; // (signal)
  /* TG68KdotC_Kernel.vhd:177:23  */
  assign lwrena = n348; // (signal)
  /* TG68KdotC_Kernel.vhd:178:16  */
  assign bwrena = n351; // (signal)
  /* TG68KdotC_Kernel.vhd:179:16  */
  assign regwrena_now = n8759; // (signal)
  /* TG68KdotC_Kernel.vhd:180:16  */
  assign rf_dest_addr = n393; // (signal)
  /* TG68KdotC_Kernel.vhd:181:16  */
  assign rf_source_addr = n431; // (signal)
  /* TG68KdotC_Kernel.vhd:182:16  */
  assign rf_source_addrd = n9332; // (signal)
  /* TG68KdotC_Kernel.vhd:184:16  */
  assign regin = n9333; // (signal)
  /* TG68KdotC_Kernel.vhd:187:16  */
  assign rdindex_a = n9337; // (signal)
  /* TG68KdotC_Kernel.vhd:188:16  */
  assign rdindex_b = n9339; // (signal)
  /* TG68KdotC_Kernel.vhd:189:16  */
  assign wr_areg = n9341; // (signal)
  /* TG68KdotC_Kernel.vhd:192:16  */
  assign addr = n994; // (signal)
  /* TG68KdotC_Kernel.vhd:193:16  */
  assign memaddr_reg = n998; // (signal)
  /* TG68KdotC_Kernel.vhd:194:16  */
  assign memaddr_delta = n993; // (signal)
  /* TG68KdotC_Kernel.vhd:195:16  */
  assign memaddr_delta_rega = n9343; // (signal)
  /* TG68KdotC_Kernel.vhd:196:16  */
  assign memaddr_delta_regb = n9345; // (signal)
  /* TG68KdotC_Kernel.vhd:197:16  */
  assign use_base = n9347; // (signal)
  /* TG68KdotC_Kernel.vhd:199:16  */
  assign ea_data = n9348; // (signal)
  /* TG68KdotC_Kernel.vhd:200:16  */
  assign op1out = n447; // (signal)
  /* TG68KdotC_Kernel.vhd:201:16  */
  assign op2out = n9349; // (signal)
  /* TG68KdotC_Kernel.vhd:202:16  */
  assign op1outbrief = n760; // (signal)
  /* TG68KdotC_Kernel.vhd:204:16  */
  assign aluout = alu_n23; // (signal)
  /* TG68KdotC_Kernel.vhd:205:16  */
  assign data_write_tmp = n9351; // (signal)
  /* TG68KdotC_Kernel.vhd:206:16  */
  assign data_write_muxin = n218; // (signal)
  /* TG68KdotC_Kernel.vhd:207:16  */
  assign data_write_mux = n227; // (signal)
  /* TG68KdotC_Kernel.vhd:208:16  */
  assign nextpass = n9352; // (signal)
  /* TG68KdotC_Kernel.vhd:209:16  */
  assign setnextpass = n8764; // (signal)
  /* TG68KdotC_Kernel.vhd:210:16  */
  assign setdispbyte = n8766; // (signal)
  /* TG68KdotC_Kernel.vhd:211:16  */
  assign setdisp = n8776; // (signal)
  /* TG68KdotC_Kernel.vhd:212:16  */
  assign regdirectsource = n7433; // (signal)
  /* TG68KdotC_Kernel.vhd:213:16  */
  assign addsub_q = alu_n22; // (signal)
  /* TG68KdotC_Kernel.vhd:214:16  */
  assign briefdata = n796; // (signal)
  /* TG68KdotC_Kernel.vhd:215:16  */
  assign c_out = alu_n21; // (signal)
  /* TG68KdotC_Kernel.vhd:218:16  */
  assign memaddr_a = n9354; // (signal)
  /* TG68KdotC_Kernel.vhd:220:16  */
  assign tg68_pc_brw = n8780; // (signal)
  /* TG68KdotC_Kernel.vhd:221:16  */
  assign tg68_pc_word = n9355; // (signal)
  /* TG68KdotC_Kernel.vhd:222:16  */
  assign getbrief = n7435; // (signal)
  /* TG68KdotC_Kernel.vhd:223:16  */
  assign brief = n9356; // (signal)
  /* TG68KdotC_Kernel.vhd:224:16  */
  assign data_is_source = n7437; // (signal)
  /* TG68KdotC_Kernel.vhd:225:16  */
  assign store_in_tmp = n9357; // (signal)
  /* TG68KdotC_Kernel.vhd:226:16  */
  assign write_back = n7823; // (signal)
  /* TG68KdotC_Kernel.vhd:227:16  */
  assign exec_write_back = n9358; // (signal)
  /* TG68KdotC_Kernel.vhd:228:16  */
  assign setstackaddr = n8794; // (signal)
  /* TG68KdotC_Kernel.vhd:229:16  */
  assign writepc = n8796; // (signal)
  /* TG68KdotC_Kernel.vhd:230:16  */
  assign writepcbig = n9359; // (signal)
  /* TG68KdotC_Kernel.vhd:231:16  */
  assign set_writepcbig = n8799; // (signal)
  /* TG68KdotC_Kernel.vhd:232:16  */
  assign writepcnext = n9360; // (signal)
  /* TG68KdotC_Kernel.vhd:233:16  */
  assign setopcode = n1122; // (signal)
  /* TG68KdotC_Kernel.vhd:234:16  */
  assign decodeopc = n9361; // (signal)
  /* TG68KdotC_Kernel.vhd:235:16  */
  assign execopc = n9362; // (signal)
  /* TG68KdotC_Kernel.vhd:236:16  */
  assign execopc_alu = n41; // (signal)
  /* TG68KdotC_Kernel.vhd:237:16  */
  assign setexecopc = n1147; // (signal)
  /* TG68KdotC_Kernel.vhd:238:16  */
  assign endopc = n9363; // (signal)
  /* TG68KdotC_Kernel.vhd:239:16  */
  assign setendopc = n1126; // (signal)
  /* TG68KdotC_Kernel.vhd:240:16  */
  assign flags = alu_n20; // (signal)
  /* TG68KdotC_Kernel.vhd:241:16  */
  assign flagssr = n9364; // (signal)
  /* TG68KdotC_Kernel.vhd:242:16  */
  assign srin = n1682; // (signal)
  /* TG68KdotC_Kernel.vhd:243:16  */
  assign exec_direct = n9365; // (signal)
  /* TG68KdotC_Kernel.vhd:244:16  */
  assign exec_tas = n9367; // (signal)
  /* TG68KdotC_Kernel.vhd:245:16  */
  assign set_exec_tas = n7447; // (signal)
  /* TG68KdotC_Kernel.vhd:247:16  */
  assign exe_condition = n9142; // (signal)
  /* TG68KdotC_Kernel.vhd:248:16  */
  assign ea_only = n7450; // (signal)
  /* TG68KdotC_Kernel.vhd:249:16  */
  assign source_areg = n8802; // (signal)
  /* TG68KdotC_Kernel.vhd:250:16  */
  assign source_lowbits = n7825; // (signal)
  /* TG68KdotC_Kernel.vhd:251:16  */
  assign source_ldrlbits = n8805; // (signal)
  /* TG68KdotC_Kernel.vhd:252:16  */
  assign source_ldrmbits = n8809; // (signal)
  /* TG68KdotC_Kernel.vhd:253:16  */
  assign source_2ndhbits = n7459; // (signal)
  /* TG68KdotC_Kernel.vhd:254:16  */
  assign source_2ndmbits = n8813; // (signal)
  /* TG68KdotC_Kernel.vhd:255:16  */
  assign source_2ndlbits = n8816; // (signal)
  /* TG68KdotC_Kernel.vhd:256:16  */
  assign dest_areg = n8821; // (signal)
  /* TG68KdotC_Kernel.vhd:257:16  */
  assign dest_ldrareg = n8823; // (signal)
  /* TG68KdotC_Kernel.vhd:258:16  */
  assign dest_ldrhbits = n8828; // (signal)
  /* TG68KdotC_Kernel.vhd:259:16  */
  assign dest_ldrlbits = n8831; // (signal)
  /* TG68KdotC_Kernel.vhd:260:16  */
  assign dest_2ndhbits = n8837; // (signal)
  /* TG68KdotC_Kernel.vhd:261:16  */
  assign dest_2ndlbits = n8841; // (signal)
  /* TG68KdotC_Kernel.vhd:262:16  */
  assign dest_hbits = n8846; // (signal)
  /* TG68KdotC_Kernel.vhd:263:16  */
  assign rot_bits = n9368; // (signal)
  /* TG68KdotC_Kernel.vhd:264:16  */
  assign set_rot_bits = n7473; // (signal)
  /* TG68KdotC_Kernel.vhd:265:16  */
  assign rot_cnt = n9369; // (signal)
  /* TG68KdotC_Kernel.vhd:266:16  */
  assign set_rot_cnt = n8848; // (signal)
  /* TG68KdotC_Kernel.vhd:267:16  */
  assign movem_actiond = n9371; // (signal)
  /* TG68KdotC_Kernel.vhd:268:16  */
  assign movem_regaddr = n9372; // (signal)
  /* TG68KdotC_Kernel.vhd:269:16  */
  assign movem_mux = n9284; // (signal)
  /* TG68KdotC_Kernel.vhd:270:16  */
  assign movem_presub = n7482; // (signal)
  /* TG68KdotC_Kernel.vhd:271:16  */
  assign movem_run = n9286; // (signal)
  /* TG68KdotC_Kernel.vhd:273:16  */
  assign set_direct_data = n8852; // (signal)
  /* TG68KdotC_Kernel.vhd:274:16  */
  assign use_direct_data = n9374; // (signal)
  /* TG68KdotC_Kernel.vhd:275:16  */
  assign direct_data = n9375; // (signal)
  /* TG68KdotC_Kernel.vhd:277:16  */
  assign set_v_flag = alu_n19; // (signal)
  /* TG68KdotC_Kernel.vhd:278:16  */
  assign set_vectoraddr = n8855; // (signal)
  /* TG68KdotC_Kernel.vhd:279:16  */
  assign writesr = n8862; // (signal)
  /* TG68KdotC_Kernel.vhd:280:16  */
  assign trap_berr = n9376; // (signal)
  /* TG68KdotC_Kernel.vhd:281:16  */
  assign trap_illegal = n8864; // (signal)
  /* TG68KdotC_Kernel.vhd:282:16  */
  assign trap_addr_error = 1'b0; // (signal)
  /* TG68KdotC_Kernel.vhd:283:16  */
  assign trap_priv = n7490; // (signal)
  /* TG68KdotC_Kernel.vhd:284:16  */
  assign trap_trace = n9377; // (signal)
  /* TG68KdotC_Kernel.vhd:285:16  */
  assign trap_1010 = n7494; // (signal)
  /* TG68KdotC_Kernel.vhd:286:16  */
  assign trap_1111 = n7497; // (signal)
  /* TG68KdotC_Kernel.vhd:287:16  */
  assign trap_trap = n7500; // (signal)
  /* TG68KdotC_Kernel.vhd:288:16  */
  assign trap_trapv = n7503; // (signal)
  /* TG68KdotC_Kernel.vhd:289:16  */
  assign trap_interrupt = n9378; // (signal)
  /* TG68KdotC_Kernel.vhd:290:16  */
  assign trapmake = n8865; // (signal)
  /* TG68KdotC_Kernel.vhd:291:16  */
  assign trapd = n9379; // (signal)
  /* TG68KdotC_Kernel.vhd:292:16  */
  assign trap_sr = n9380; // (signal)
  /* TG68KdotC_Kernel.vhd:293:16  */
  assign make_trace = n9381; // (signal)
  /* TG68KdotC_Kernel.vhd:294:16  */
  assign make_berr = n9382; // (signal)
  /* TG68KdotC_Kernel.vhd:295:16  */
  assign usestackframe2 = n9383; // (signal)
  /* TG68KdotC_Kernel.vhd:297:16  */
  assign set_stop = n7512; // (signal)
  /* TG68KdotC_Kernel.vhd:298:16  */
  assign stop = n9384; // (signal)
  /* TG68KdotC_Kernel.vhd:299:16  */
  assign trap_vector = n9386; // (signal)
  /* TG68KdotC_Kernel.vhd:300:16  */
  assign trap_vector_vbr = n838; // (signal)
  /* TG68KdotC_Kernel.vhd:301:16  */
  assign usp = n9388; // (signal)
  /* TG68KdotC_Kernel.vhd:306:16  */
  assign ipl_nr = n1149; // (signal)
  /* TG68KdotC_Kernel.vhd:307:16  */
  assign ripl_nr = n9389; // (signal)
  /* TG68KdotC_Kernel.vhd:308:16  */
  assign ipl_vec = n9390; // (signal)
  /* TG68KdotC_Kernel.vhd:309:16  */
  assign interrupt = n9391; // (signal)
  /* TG68KdotC_Kernel.vhd:310:16  */
  assign setinterrupt = n1129; // (signal)
  /* TG68KdotC_Kernel.vhd:311:16  */
  assign svmode = n9392; // (signal)
  /* TG68KdotC_Kernel.vhd:312:16  */
  assign presvmode = n9393; // (signal)
  /* TG68KdotC_Kernel.vhd:313:16  */
  assign suppress_base = n9394; // (signal)
  /* TG68KdotC_Kernel.vhd:314:16  */
  assign set_suppress_base = n8868; // (signal)
  /* TG68KdotC_Kernel.vhd:315:16  */
  assign set_z_error = n8870; // (signal)
  /* TG68KdotC_Kernel.vhd:316:16  */
  assign z_error = n9395; // (signal)
  /* TG68KdotC_Kernel.vhd:317:16  */
  assign ea_build_now = n7789; // (signal)
  /* TG68KdotC_Kernel.vhd:318:16  */
  assign build_logical = n7518; // (signal)
  /* TG68KdotC_Kernel.vhd:319:16  */
  assign build_bcd = n7521; // (signal)
  /* TG68KdotC_Kernel.vhd:321:16  */
  assign data_read = n9396; // (signal)
  /* TG68KdotC_Kernel.vhd:322:16  */
  assign bf_ext_in = n9398; // (signal)
  /* TG68KdotC_Kernel.vhd:323:16  */
  assign bf_ext_out = alu_n17; // (signal)
  /* TG68KdotC_Kernel.vhd:325:16  */
  assign long_start = n211; // (signal)
  /* TG68KdotC_Kernel.vhd:326:16  */
  assign long_start_alu = n39; // (signal)
  /* TG68KdotC_Kernel.vhd:327:16  */
  assign non_aligned = n53; // (signal)
  /* TG68KdotC_Kernel.vhd:328:16  */
  assign check_aligned = n7524; // (signal)
  /* TG68KdotC_Kernel.vhd:329:16  */
  assign long_done = n213; // (signal)
  /* TG68KdotC_Kernel.vhd:330:16  */
  assign memmask = n9399; // (signal)
  /* TG68KdotC_Kernel.vhd:331:16  */
  assign set_memmask = n1666; // (signal)
  /* TG68KdotC_Kernel.vhd:332:16  */
  assign memread = n9400; // (signal)
  /* TG68KdotC_Kernel.vhd:333:16  */
  assign wbmemmask = n9401; // (signal)
  /* TG68KdotC_Kernel.vhd:334:16  */
  assign memmaskmux = n66; // (signal)
  /* TG68KdotC_Kernel.vhd:335:16  */
  assign oddout = n9402; // (signal)
  /* TG68KdotC_Kernel.vhd:336:16  */
  assign set_oddout = n1601; // (signal)
  /* TG68KdotC_Kernel.vhd:337:16  */
  assign pcbase = n9403; // (signal)
  /* TG68KdotC_Kernel.vhd:338:16  */
  assign set_pcbase = n2037; // (signal)
  /* TG68KdotC_Kernel.vhd:340:16  */
  assign last_data_read = n9404; // (signal)
  /* TG68KdotC_Kernel.vhd:341:16  */
  assign last_data_in = n9405; // (signal)
  /* TG68KdotC_Kernel.vhd:343:16  */
  assign bf_offset = n9406; // (signal)
  /* TG68KdotC_Kernel.vhd:344:16  */
  assign bf_width = n9407; // (signal)
  /* TG68KdotC_Kernel.vhd:345:16  */
  assign bf_bhits = n1599; // (signal)
  /* TG68KdotC_Kernel.vhd:346:16  */
  assign bf_shift = n1646; // (signal)
  /* TG68KdotC_Kernel.vhd:347:16  */
  assign alu_width = n9408; // (signal)
  /* TG68KdotC_Kernel.vhd:348:16  */
  assign alu_bf_shift = n9409; // (signal)
  /* TG68KdotC_Kernel.vhd:349:16  */
  assign bf_loffset = n9410; // (signal)
  /* TG68KdotC_Kernel.vhd:350:16  */
  assign bf_full_offset = n1589; // (signal)
  /* TG68KdotC_Kernel.vhd:351:16  */
  assign alu_bf_ffo_offset = n9411; // (signal)
  /* TG68KdotC_Kernel.vhd:352:16  */
  assign alu_bf_loffset = n9412; // (signal)
  /* TG68KdotC_Kernel.vhd:354:16  */
  assign movec_data = n9037; // (signal)
  /* TG68KdotC_Kernel.vhd:355:16  */
  assign vbr = n9413; // (signal)
  /* TG68KdotC_Kernel.vhd:356:16  */
  assign cacr = n9414; // (signal)
  /* TG68KdotC_Kernel.vhd:357:16  */
  assign dfc = n9415; // (signal)
  /* TG68KdotC_Kernel.vhd:358:16  */
  assign sfc = n9416; // (signal)
  /* TG68KdotC_Kernel.vhd:361:16  */
  assign set = n9417; // (signal)
  /* TG68KdotC_Kernel.vhd:362:16  */
  assign set_exec = n9418; // (signal)
  /* TG68KdotC_Kernel.vhd:363:16  */
  assign exec = n9420; // (signal)
  /* TG68KdotC_Kernel.vhd:365:16  */
  assign micro_state = n9421; // (signal)
  /* TG68KdotC_Kernel.vhd:366:16  */
  assign next_micro_state = n8971; // (signal)
  /* TG68KdotC_Kernel.vhd:405:49  */
  assign n15 = last_data_read[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:406:39  */
  assign n16 = data_read[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:414:45  */
  assign n18 = alu_bf_loffset[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:372:1  */
  tg68k_alu_2_1_2_2 alu (
    .clk(clk),
    .reset(reset),
    .clkena_lw(clkena_lw),
    .cpu(CPU),
    .execopc(execopc_alu),
    .decodeopc(decodeopc),
    .exe_condition(exe_condition),
    .exec_tas(exec_tas),
    .long_start(long_start_alu),
    .non_aligned(non_aligned),
    .check_aligned(check_aligned),
    .movem_presub(movem_presub),
    .set_stop(set_stop),
    .z_error(z_error),
    .rot_bits(rot_bits),
    .exec(exec),
    .op1out(op1out),
    .op2out(op2out),
    .reg_qa(reg_qa),
    .reg_qb(reg_qb),
    .opcode(opcode),
    .exe_opcode(exe_opcode),
    .exe_datatype(exe_datatype),
    .sndopc(sndopc),
    .last_data_read(n15),
    .data_read(n16),
    .flagssr(flagssr),
    .micro_state(micro_state),
    .bf_ext_in(bf_ext_in),
    .bf_shift(alu_bf_shift),
    .bf_width(alu_width),
    .bf_ffo_offset(alu_bf_ffo_offset),
    .bf_loffset(n18),
    .bf_ext_out(alu_n17),
    .set_v_flag(alu_n19),
    .flags(alu_n20),
    .c_out(alu_n21),
    .addsub_q(alu_n22),
    .aluout(alu_n23));
  /* TG68KdotC_Kernel.vhd:424:35  */
  assign n36 = memmaskmux[3]; // extract
  /* TG68KdotC_Kernel.vhd:424:21  */
  assign n37 = ~n36;
  /* TG68KdotC_Kernel.vhd:426:48  */
  assign n38 = memmaskmux[3]; // extract
  /* TG68KdotC_Kernel.vhd:426:34  */
  assign n39 = ~n38;
  /* TG68KdotC_Kernel.vhd:427:39  */
  assign n40 = exec[84]; // extract
  /* TG68KdotC_Kernel.vhd:427:32  */
  assign n41 = execopc | n40;
  /* TG68KdotC_Kernel.vhd:431:31  */
  assign n44 = memmaskmux[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:431:44  */
  assign n46 = n44 == 2'b01;
  /* TG68KdotC_Kernel.vhd:431:66  */
  assign n47 = memmaskmux[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:431:79  */
  assign n49 = n47 == 2'b10;
  /* TG68KdotC_Kernel.vhd:431:52  */
  assign n50 = n46 | n49;
  /* TG68KdotC_Kernel.vhd:431:17  */
  assign n53 = n50 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:441:30  */
  assign n58 = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:441:20  */
  assign n59 = n58 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:443:35  */
  assign n62 = exec[74]; // extract
  /* TG68KdotC_Kernel.vhd:443:26  */
  assign n63 = n62 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:447:40  */
  assign n65 = addr[0]; // extract
  /* TG68KdotC_Kernel.vhd:447:31  */
  assign n66 = n65 ? memmask : n69;
  /* TG68KdotC_Kernel.vhd:447:62  */
  assign n67 = memmask[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:447:75  */
  assign n69 = {n67, 1'b1};
  /* TG68KdotC_Kernel.vhd:448:27  */
  assign n70 = memmaskmux[5]; // extract
  /* TG68KdotC_Kernel.vhd:449:27  */
  assign n71 = memmaskmux[4]; // extract
  /* TG68KdotC_Kernel.vhd:450:59  */
  assign n73 = memmaskmux[3]; // extract
  /* TG68KdotC_Kernel.vhd:450:45  */
  assign n74 = n73 & clkena_in;
  /* TG68KdotC_Kernel.vhd:450:26  */
  assign n75 = n74 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:451:44  */
  assign n78 = trap_berr & setopcode;
  /* TG68KdotC_Kernel.vhd:451:25  */
  assign n79 = n78 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:455:26  */
  assign n83 = ~nReset;
  /* TG68KdotC_Kernel.vhd:460:55  */
  assign n85 = syncreset[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:460:67  */
  assign n87 = {n85, 1'b1};
  /* TG68KdotC_Kernel.vhd:461:55  */
  assign n88 = syncreset[3]; // extract
  /* TG68KdotC_Kernel.vhd:461:42  */
  assign n89 = ~n88;
  /* TG68KdotC_Kernel.vhd:465:52  */
  assign n99 = CPU[0]; // extract
  /* TG68KdotC_Kernel.vhd:465:60  */
  assign n101 = 1'b1 & n99;
  /* TG68KdotC_Kernel.vhd:465:45  */
  assign n103 = 1'b0 | n101;
  /* TG68KdotC_Kernel.vhd:465:25  */
  assign n106 = n103 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:475:30  */
  assign n111 = memmaskmux[4]; // extract
  /* TG68KdotC_Kernel.vhd:475:33  */
  assign n112 = ~n111;
  /* TG68KdotC_Kernel.vhd:476:50  */
  assign n113 = last_data_in[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:476:63  */
  assign n114 = {n113, data_in};
  /* TG68KdotC_Kernel.vhd:478:50  */
  assign n115 = last_data_in[23:0]; // extract
  /* TG68KdotC_Kernel.vhd:478:71  */
  assign n116 = data_in[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:478:63  */
  assign n117 = {n115, n116};
  /* TG68KdotC_Kernel.vhd:475:17  */
  assign n118 = n112 ? n114 : n117;
  /* TG68KdotC_Kernel.vhd:480:27  */
  assign n119 = memread[0]; // extract
  /* TG68KdotC_Kernel.vhd:480:46  */
  assign n120 = memread[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:480:58  */
  assign n122 = n120 == 2'b10;
  /* TG68KdotC_Kernel.vhd:480:78  */
  assign n123 = memmaskmux[4]; // extract
  /* TG68KdotC_Kernel.vhd:480:64  */
  assign n124 = n123 & n122;
  /* TG68KdotC_Kernel.vhd:480:35  */
  assign n125 = n119 | n124;
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n126 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n127 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n128 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n129 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n130 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n131 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n132 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n133 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n134 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n135 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n136 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n137 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n138 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n139 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n140 = data_read[15]; // extract
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n141 = data_read[15]; // extract
  assign n142 = {n126, n127, n128, n129};
  assign n143 = {n130, n131, n132, n133};
  assign n144 = {n134, n135, n136, n137};
  assign n145 = {n138, n139, n140, n141};
  assign n146 = {n142, n143, n144, n145};
  assign n147 = n118[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:480:17  */
  assign n148 = n125 ? n146 : n147;
  assign n149 = n118[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:485:51  */
  assign n152 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:485:42  */
  assign n153 = n152 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:486:46  */
  assign n154 = memmaskmux[4]; // extract
  /* TG68KdotC_Kernel.vhd:486:49  */
  assign n155 = ~n154;
  /* TG68KdotC_Kernel.vhd:487:66  */
  assign n156 = last_data_in[23:16]; // extract
  /* TG68KdotC_Kernel.vhd:489:66  */
  assign n157 = last_data_in[31:24]; // extract
  /* TG68KdotC_Kernel.vhd:486:33  */
  assign n158 = n155 ? n156 : n157;
  /* TG68KdotC_Kernel.vhd:495:41  */
  assign n161 = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:495:54  */
  assign n162 = exec[38]; // extract
  /* TG68KdotC_Kernel.vhd:495:47  */
  assign n163 = n161 | n162;
  /* TG68KdotC_Kernel.vhd:497:49  */
  assign n164 = state[1]; // extract
  /* TG68KdotC_Kernel.vhd:497:52  */
  assign n165 = ~n164;
  /* TG68KdotC_Kernel.vhd:497:68  */
  assign n166 = memmask[1]; // extract
  /* TG68KdotC_Kernel.vhd:497:71  */
  assign n167 = ~n166;
  /* TG68KdotC_Kernel.vhd:497:57  */
  assign n168 = n167 & n165;
  /* TG68KdotC_Kernel.vhd:499:52  */
  assign n169 = state[1]; // extract
  /* TG68KdotC_Kernel.vhd:499:55  */
  assign n170 = ~n169;
  /* TG68KdotC_Kernel.vhd:499:70  */
  assign n171 = memread[1]; // extract
  /* TG68KdotC_Kernel.vhd:499:60  */
  assign n172 = n170 | n171;
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n173 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n174 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n175 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n176 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n177 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n178 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n179 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n180 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n181 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n182 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n183 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n184 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n185 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n186 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n187 = data_in[15]; // extract
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n188 = data_in[15]; // extract
  assign n189 = {n173, n174, n175, n176};
  assign n190 = {n177, n178, n179, n180};
  assign n191 = {n181, n182, n183, n184};
  assign n192 = {n185, n186, n187, n188};
  assign n193 = {n189, n190, n191, n192};
  assign n194 = data_read[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:499:41  */
  assign n195 = n172 ? n193 : n194;
  /* TG68KdotC_Kernel.vhd:497:41  */
  assign n196 = n168 ? last_opc_read : n195;
  assign n197 = data_read[15:0]; // extract
  assign n198 = {n196, n197};
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n199 = n202 ? n198 : last_data_read;
  /* TG68KdotC_Kernel.vhd:503:61  */
  assign n200 = last_data_in[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:503:74  */
  assign n201 = {n200, data_in};
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n202 = n163 & clkena_in;
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n203 = clkena_in ? n201 : last_data_in;
  /* TG68KdotC_Kernel.vhd:492:25  */
  assign n205 = reset ? 32'b00000000000000000000000000000000 : n199;
  /* TG68KdotC_Kernel.vhd:492:25  */
  assign n206 = reset ? last_data_in : n203;
  /* TG68KdotC_Kernel.vhd:507:65  */
  assign n210 = memmask[1]; // extract
  /* TG68KdotC_Kernel.vhd:507:54  */
  assign n211 = ~n210;
  /* TG68KdotC_Kernel.vhd:508:64  */
  assign n212 = memread[1]; // extract
  /* TG68KdotC_Kernel.vhd:508:53  */
  assign n213 = ~n212;
  /* TG68KdotC_Kernel.vhd:514:24  */
  assign n217 = exec[40]; // extract
  /* TG68KdotC_Kernel.vhd:514:17  */
  assign n218 = n217 ? reg_qb : data_write_tmp;
  /* TG68KdotC_Kernel.vhd:527:39  */
  assign n219 = addr[0]; // extract
  /* TG68KdotC_Kernel.vhd:527:34  */
  assign n220 = oddout == n219;
  /* TG68KdotC_Kernel.vhd:528:61  */
  assign n222 = {8'bX, bf_ext_out};
  /* TG68KdotC_Kernel.vhd:528:72  */
  assign n223 = {n222, data_write_muxin};
  /* TG68KdotC_Kernel.vhd:530:61  */
  assign n224 = {bf_ext_out, data_write_muxin};
  /* TG68KdotC_Kernel.vhd:530:78  */
  assign n226 = {n224, 8'bX};
  /* TG68KdotC_Kernel.vhd:527:25  */
  assign n227 = n220 ? n223 : n226;
  /* TG68KdotC_Kernel.vhd:534:30  */
  assign n228 = memmaskmux[1]; // extract
  /* TG68KdotC_Kernel.vhd:534:33  */
  assign n229 = ~n228;
  /* TG68KdotC_Kernel.vhd:535:53  */
  assign n230 = data_write_mux[47:32]; // extract
  /* TG68KdotC_Kernel.vhd:536:33  */
  assign n231 = memmaskmux[3]; // extract
  /* TG68KdotC_Kernel.vhd:536:36  */
  assign n232 = ~n231;
  /* TG68KdotC_Kernel.vhd:537:53  */
  assign n233 = data_write_mux[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:540:38  */
  assign n234 = memmaskmux[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:540:51  */
  assign n236 = n234 == 2'b10;
  /* TG68KdotC_Kernel.vhd:541:61  */
  assign n237 = data_write_mux[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:541:90  */
  assign n238 = data_write_mux[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:541:74  */
  assign n239 = {n237, n238};
  /* TG68KdotC_Kernel.vhd:542:41  */
  assign n240 = memmaskmux[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:542:54  */
  assign n242 = n240 == 2'b01;
  /* TG68KdotC_Kernel.vhd:543:61  */
  assign n243 = data_write_mux[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:543:91  */
  assign n244 = data_write_mux[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:543:75  */
  assign n245 = {n243, n244};
  /* TG68KdotC_Kernel.vhd:545:61  */
  assign n246 = data_write_mux[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:542:25  */
  assign n247 = n242 ? n245 : n246;
  /* TG68KdotC_Kernel.vhd:540:25  */
  assign n248 = n236 ? n239 : n247;
  /* TG68KdotC_Kernel.vhd:536:17  */
  assign n249 = n232 ? n233 : n248;
  /* TG68KdotC_Kernel.vhd:534:17  */
  assign n250 = n229 ? n230 : n249;
  /* TG68KdotC_Kernel.vhd:548:24  */
  assign n251 = exec[72]; // extract
  /* TG68KdotC_Kernel.vhd:549:65  */
  assign n252 = data_write_tmp[15:8]; // extract
  assign n253 = n250[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:548:17  */
  assign n254 = n251 ? n252 : n253;
  assign n255 = n250[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:563:56  */
  assign n268 = rf_dest_addr[3]; // extract
  /* TG68KdotC_Kernel.vhd:570:40  */
  assign n276 = exec[65]; // extract
  /* TG68KdotC_Kernel.vhd:561:21  */
  assign n279 = wwrena & clkena_lw;
  /* TG68KdotC_Kernel.vhd:561:21  */
  assign n283 = n276 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:583:24  */
  assign n293 = exec[30]; // extract
  /* TG68KdotC_Kernel.vhd:585:27  */
  assign n294 = exec[62]; // extract
  /* TG68KdotC_Kernel.vhd:585:44  */
  assign n295 = ea_only & n294;
  /* TG68KdotC_Kernel.vhd:587:27  */
  assign n296 = exec[66]; // extract
  /* TG68KdotC_Kernel.vhd:589:27  */
  assign n297 = exec[32]; // extract
  /* TG68KdotC_Kernel.vhd:589:17  */
  assign n298 = n297 ? movec_data : aluout;
  /* TG68KdotC_Kernel.vhd:587:17  */
  assign n299 = n296 ? usp : n298;
  /* TG68KdotC_Kernel.vhd:585:17  */
  assign n300 = n295 ? memaddr_a : n299;
  /* TG68KdotC_Kernel.vhd:583:17  */
  assign n301 = n293 ? memaddr : n300;
  /* TG68KdotC_Kernel.vhd:594:53  */
  assign n302 = reg_qa[15:8]; // extract
  assign n303 = n301[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:593:17  */
  assign n304 = bwrena ? n302 : n303;
  assign n305 = n301[31:16]; // extract
  assign n306 = n301[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:596:26  */
  assign n307 = ~lwrena;
  /* TG68KdotC_Kernel.vhd:597:54  */
  assign n308 = reg_qa[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:596:17  */
  assign n309 = n307 ? n308 : n305;
  /* TG68KdotC_Kernel.vhd:603:24  */
  assign n310 = exec[47]; // extract
  /* TG68KdotC_Kernel.vhd:603:44  */
  assign n311 = exec[46]; // extract
  /* TG68KdotC_Kernel.vhd:603:37  */
  assign n312 = n310 | n311;
  /* TG68KdotC_Kernel.vhd:603:65  */
  assign n313 = exec[41]; // extract
  /* TG68KdotC_Kernel.vhd:603:58  */
  assign n314 = n312 | n313;
  /* TG68KdotC_Kernel.vhd:608:27  */
  assign n315 = exec[34]; // extract
  /* TG68KdotC_Kernel.vhd:611:33  */
  assign n317 = exe_datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:614:56  */
  assign n318 = wr_areg | movem_actiond;
  /* TG68KdotC_Kernel.vhd:614:41  */
  assign n321 = n318 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:613:33  */
  assign n323 = exe_datatype == 2'b01;
  assign n324 = {n323, n317};
  /* TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n324)
      2'b10: n327 = n321;
      2'b01: n327 = 1'b0;
      default: n327 = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n324)
      2'b10: n330 = 1'b0;
      2'b01: n330 = 1'b1;
      default: n330 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n333 = n315 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n335 = n315 ? n327 : 1'b0;
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n337 = n315 ? n330 : 1'b0;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n339 = regwrena_now ? 1'b1 : n333;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n341 = regwrena_now ? 1'b0 : n335;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n343 = regwrena_now ? 1'b0 : n337;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n345 = n314 ? 1'b1 : n339;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n348 = n314 ? 1'b1 : n341;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n351 = n314 ? 1'b0 : n343;
  /* TG68KdotC_Kernel.vhd:628:24  */
  assign n356 = exec[69]; // extract
  /* TG68KdotC_Kernel.vhd:630:26  */
  assign n357 = set[70]; // extract
  /* TG68KdotC_Kernel.vhd:631:46  */
  assign n358 = brief[15:12]; // extract
  /* TG68KdotC_Kernel.vhd:632:26  */
  assign n359 = set[29]; // extract
  /* TG68KdotC_Kernel.vhd:634:59  */
  assign n360 = sndopc[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:634:52  */
  assign n362 = {1'b0, n360};
  /* TG68KdotC_Kernel.vhd:639:60  */
  assign n363 = sndopc[14:12]; // extract
  /* TG68KdotC_Kernel.vhd:639:53  */
  assign n364 = {dest_ldrareg, n363};
  /* TG68KdotC_Kernel.vhd:641:55  */
  assign n365 = last_data_read[15:12]; // extract
  /* TG68KdotC_Kernel.vhd:643:59  */
  assign n366 = last_data_read[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:643:44  */
  assign n368 = {1'b0, n366};
  /* TG68KdotC_Kernel.vhd:645:51  */
  assign n369 = sndopc[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:645:44  */
  assign n371 = {1'b0, n369};
  /* TG68KdotC_Kernel.vhd:649:57  */
  assign n372 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:649:50  */
  assign n373 = {dest_areg, n372};
  /* TG68KdotC_Kernel.vhd:651:34  */
  assign n374 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:651:46  */
  assign n376 = n374 == 3'b000;
  /* TG68KdotC_Kernel.vhd:651:53  */
  assign n377 = n376 | data_is_source;
  /* TG68KdotC_Kernel.vhd:652:65  */
  assign n378 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:652:58  */
  assign n379 = {dest_areg, n378};
  /* TG68KdotC_Kernel.vhd:654:59  */
  assign n380 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:654:52  */
  assign n382 = {1'b1, n380};
  /* TG68KdotC_Kernel.vhd:651:25  */
  assign n383 = n377 ? n379 : n382;
  /* TG68KdotC_Kernel.vhd:648:17  */
  assign n384 = dest_hbits ? n373 : n383;
  /* TG68KdotC_Kernel.vhd:646:17  */
  assign n386 = setstackaddr ? 4'b1111 : n384;
  /* TG68KdotC_Kernel.vhd:644:17  */
  assign n387 = dest_2ndlbits ? n371 : n386;
  /* TG68KdotC_Kernel.vhd:642:17  */
  assign n388 = dest_ldrlbits ? n368 : n387;
  /* TG68KdotC_Kernel.vhd:640:17  */
  assign n389 = dest_ldrhbits ? n365 : n388;
  /* TG68KdotC_Kernel.vhd:638:17  */
  assign n390 = dest_2ndhbits ? n364 : n389;
  /* TG68KdotC_Kernel.vhd:632:17  */
  assign n391 = n359 ? n362 : n390;
  /* TG68KdotC_Kernel.vhd:630:17  */
  assign n392 = n357 ? n358 : n391;
  /* TG68KdotC_Kernel.vhd:628:17  */
  assign n393 = n356 ? rf_source_addrd : n392;
  /* TG68KdotC_Kernel.vhd:664:24  */
  assign n397 = exec[69]; // extract
  /* TG68KdotC_Kernel.vhd:664:49  */
  assign n398 = set[69]; // extract
  /* TG68KdotC_Kernel.vhd:664:43  */
  assign n399 = n397 | n398;
  /* TG68KdotC_Kernel.vhd:666:65  */
  assign n401 = movem_regaddr ^ 4'b1111;
  /* TG68KdotC_Kernel.vhd:665:25  */
  assign n402 = movem_presub ? n401 : movem_regaddr;
  /* TG68KdotC_Kernel.vhd:671:53  */
  assign n403 = sndopc[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:671:46  */
  assign n405 = {1'b0, n403};
  /* TG68KdotC_Kernel.vhd:673:53  */
  assign n406 = sndopc[14:12]; // extract
  /* TG68KdotC_Kernel.vhd:673:46  */
  assign n408 = {1'b0, n406};
  /* TG68KdotC_Kernel.vhd:675:53  */
  assign n409 = sndopc[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:675:46  */
  assign n411 = {1'b0, n409};
  /* TG68KdotC_Kernel.vhd:677:61  */
  assign n412 = last_data_read[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:677:46  */
  assign n414 = {1'b0, n412};
  /* TG68KdotC_Kernel.vhd:679:61  */
  assign n415 = last_data_read[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:679:46  */
  assign n417 = {1'b0, n415};
  /* TG68KdotC_Kernel.vhd:681:61  */
  assign n418 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:681:54  */
  assign n419 = {source_areg, n418};
  /* TG68KdotC_Kernel.vhd:682:27  */
  assign n420 = exec[36]; // extract
  /* TG68KdotC_Kernel.vhd:685:61  */
  assign n421 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:685:54  */
  assign n422 = {source_areg, n421};
  /* TG68KdotC_Kernel.vhd:682:17  */
  assign n424 = n420 ? 4'b1111 : n422;
  /* TG68KdotC_Kernel.vhd:680:17  */
  assign n425 = source_lowbits ? n419 : n424;
  /* TG68KdotC_Kernel.vhd:678:17  */
  assign n426 = source_ldrmbits ? n417 : n425;
  /* TG68KdotC_Kernel.vhd:676:17  */
  assign n427 = source_ldrlbits ? n414 : n426;
  /* TG68KdotC_Kernel.vhd:674:17  */
  assign n428 = source_2ndmbits ? n411 : n427;
  /* TG68KdotC_Kernel.vhd:672:17  */
  assign n429 = source_2ndhbits ? n408 : n428;
  /* TG68KdotC_Kernel.vhd:670:17  */
  assign n430 = source_2ndlbits ? n405 : n429;
  /* TG68KdotC_Kernel.vhd:664:17  */
  assign n431 = n399 ? n402 : n430;
  /* TG68KdotC_Kernel.vhd:695:24  */
  assign n435 = exec[54]; // extract
  /* TG68KdotC_Kernel.vhd:697:27  */
  assign n436 = exec[26]; // extract
  /* TG68KdotC_Kernel.vhd:697:45  */
  assign n437 = store_in_tmp & n436;
  /* TG68KdotC_Kernel.vhd:699:27  */
  assign n438 = exec[69]; // extract
  /* TG68KdotC_Kernel.vhd:699:59  */
  assign n439 = memmaskmux[3]; // extract
  /* TG68KdotC_Kernel.vhd:699:62  */
  assign n440 = ~n439;
  /* TG68KdotC_Kernel.vhd:699:46  */
  assign n441 = n438 | n440;
  /* TG68KdotC_Kernel.vhd:699:74  */
  assign n442 = exec[39]; // extract
  /* TG68KdotC_Kernel.vhd:699:67  */
  assign n443 = n441 | n442;
  /* TG68KdotC_Kernel.vhd:699:17  */
  assign n444 = n443 ? addr : reg_qa;
  /* TG68KdotC_Kernel.vhd:697:17  */
  assign n445 = n437 ? ea_data : n444;
  /* TG68KdotC_Kernel.vhd:695:17  */
  assign n447 = n435 ? 32'b00000000000000000000000000000000 : n445;
  /* TG68KdotC_Kernel.vhd:710:46  */
  assign n451 = reg_qb[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n452 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n453 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n454 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n455 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n456 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n457 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n458 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n459 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n460 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n461 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n462 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n463 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n464 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n465 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n466 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n467 = op2out[15]; // extract
  assign n468 = {n452, n453, n454, n455};
  assign n469 = {n456, n457, n458, n459};
  assign n470 = {n460, n461, n462, n463};
  assign n471 = {n464, n465, n466, n467};
  assign n472 = {n468, n469, n470, n471};
  /* TG68KdotC_Kernel.vhd:712:24  */
  assign n473 = exec[53]; // extract
  /* TG68KdotC_Kernel.vhd:714:51  */
  assign n475 = exec[61]; // extract
  /* TG68KdotC_Kernel.vhd:714:61  */
  assign n476 = execopc & n475;
  /* TG68KdotC_Kernel.vhd:714:43  */
  assign n477 = use_direct_data | n476;
  /* TG68KdotC_Kernel.vhd:714:85  */
  assign n478 = exec[29]; // extract
  /* TG68KdotC_Kernel.vhd:714:78  */
  assign n479 = n477 | n478;
  /* TG68KdotC_Kernel.vhd:716:28  */
  assign n480 = exec[26]; // extract
  /* TG68KdotC_Kernel.vhd:716:41  */
  assign n481 = ~n480;
  /* TG68KdotC_Kernel.vhd:716:46  */
  assign n482 = store_in_tmp & n481;
  /* TG68KdotC_Kernel.vhd:716:75  */
  assign n483 = exec[27]; // extract
  /* TG68KdotC_Kernel.vhd:716:68  */
  assign n484 = n482 | n483;
  /* TG68KdotC_Kernel.vhd:718:27  */
  assign n485 = exec[1]; // extract
  /* TG68KdotC_Kernel.vhd:719:57  */
  assign n486 = exe_opcode[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n487 = exe_opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n488 = exe_opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n489 = exe_opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n490 = exe_opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n491 = exe_opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n492 = exe_opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n493 = exe_opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n494 = exe_opcode[7]; // extract
  assign n495 = {n487, n488, n489, n490};
  assign n496 = {n491, n492, n493, n494};
  assign n497 = {n495, n496};
  /* TG68KdotC_Kernel.vhd:721:27  */
  assign n498 = exec[4]; // extract
  /* TG68KdotC_Kernel.vhd:722:57  */
  assign n499 = exe_opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:723:38  */
  assign n500 = exe_opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:723:51  */
  assign n502 = n500 == 3'b000;
  /* TG68KdotC_Kernel.vhd:723:25  */
  assign n505 = n502 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:729:35  */
  assign n508 = exe_datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:729:49  */
  assign n509 = exec[11]; // extract
  /* TG68KdotC_Kernel.vhd:729:57  */
  assign n510 = ~n509;
  /* TG68KdotC_Kernel.vhd:729:41  */
  assign n511 = n510 & n508;
  /* TG68KdotC_Kernel.vhd:730:55  */
  assign n512 = reg_qb[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:729:17  */
  assign n513 = n511 ? n512 : n472;
  assign n514 = {12'b000000000000, n505, n499};
  /* TG68KdotC_Kernel.vhd:721:17  */
  assign n515 = n498 ? n514 : n451;
  /* TG68KdotC_Kernel.vhd:721:17  */
  assign n516 = n498 ? n472 : n513;
  assign n517 = {n516, n515};
  assign n518 = {n497, n486};
  assign n519 = n517[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:718:17  */
  assign n520 = n485 ? n518 : n519;
  assign n521 = n517[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:718:17  */
  assign n522 = n485 ? n472 : n521;
  assign n523 = {n522, n520};
  /* TG68KdotC_Kernel.vhd:716:17  */
  assign n524 = n484 ? ea_data : n523;
  /* TG68KdotC_Kernel.vhd:714:17  */
  assign n525 = n479 ? data_write_tmp : n524;
  assign n526 = n525[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n527 = n473 ? 16'b1111111111111111 : n526;
  assign n528 = n525[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n529 = n473 ? n472 : n528;
  /* TG68KdotC_Kernel.vhd:732:24  */
  assign n530 = exec[88]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n531 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n532 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n533 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n534 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n535 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n536 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n537 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n538 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n539 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n540 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n541 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n542 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n543 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n544 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n545 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n546 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n547 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n548 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n549 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n550 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n551 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n552 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n553 = op2out[7]; // extract
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n554 = op2out[7]; // extract
  assign n555 = {n531, n532, n533, n534};
  assign n556 = {n535, n536, n537, n538};
  assign n557 = {n539, n540, n541, n542};
  assign n558 = {n543, n544, n545, n546};
  assign n559 = {n547, n548, n549, n550};
  assign n560 = {n551, n552, n553, n554};
  assign n561 = {n555, n556, n557, n558};
  assign n562 = {n559, n560};
  assign n563 = {n561, n562};
  assign n564 = n527[15:8]; // extract
  assign n565 = {n529, n564};
  /* TG68KdotC_Kernel.vhd:732:17  */
  assign n566 = n530 ? n563 : n565;
  assign n567 = n527[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:753:40  */
  assign n572 = exec[82]; // extract
  /* TG68KdotC_Kernel.vhd:753:33  */
  assign n574 = n572 ? 1'b1 : use_direct_data;
  /* TG68KdotC_Kernel.vhd:759:56  */
  assign n575 = set[27]; // extract
  /* TG68KdotC_Kernel.vhd:759:50  */
  assign n576 = endopc | n575;
  /* TG68KdotC_Kernel.vhd:759:33  */
  assign n578 = n576 ? 1'b0 : n574;
  /* TG68KdotC_Kernel.vhd:756:33  */
  assign n580 = set_direct_data ? 1'b1 : n578;
  /* TG68KdotC_Kernel.vhd:756:33  */
  assign n583 = set_direct_data ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:762:56  */
  assign n585 = set_exec[0]; // extract
  /* TG68KdotC_Kernel.vhd:769:41  */
  assign n587 = set_z_error ? 1'b1 : z_error;
  /* TG68KdotC_Kernel.vhd:772:52  */
  assign n588 = set_exec[0]; // extract
  /* TG68KdotC_Kernel.vhd:772:75  */
  assign n590 = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:772:66  */
  assign n591 = n590 & n588;
  /* TG68KdotC_Kernel.vhd:772:41  */
  assign n593 = n591 ? 1'b1 : n580;
  /* TG68KdotC_Kernel.vhd:776:49  */
  assign n595 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:776:62  */
  assign n596 = exec[80]; // extract
  /* TG68KdotC_Kernel.vhd:776:55  */
  assign n597 = n595 | n596;
  /* TG68KdotC_Kernel.vhd:776:41  */
  assign n599 = n597 ? 1'b1 : store_in_tmp;
  /* TG68KdotC_Kernel.vhd:779:69  */
  assign n601 = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:779:60  */
  assign n602 = n601 & direct_data;
  /* TG68KdotC_Kernel.vhd:779:41  */
  assign n604 = n602 ? 1'b1 : n599;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n606 = endopc ? 1'b0 : n604;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n608 = endopc ? 1'b0 : writepcnext;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n609 = endopc ? n580 : n593;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n611 = endopc ? 1'b0 : n587;
  /* TG68KdotC_Kernel.vhd:784:41  */
  assign n613 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:784:55  */
  assign n614 = exec[79]; // extract
  /* TG68KdotC_Kernel.vhd:784:69  */
  assign n615 = ~n614;
  /* TG68KdotC_Kernel.vhd:784:47  */
  assign n616 = n615 & n613;
  /* TG68KdotC_Kernel.vhd:786:43  */
  assign n617 = exec[71]; // extract
  /* TG68KdotC_Kernel.vhd:788:43  */
  assign n618 = exec[44]; // extract
  /* TG68KdotC_Kernel.vhd:788:92  */
  assign n620 = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:788:83  */
  assign n621 = n620 & direct_data;
  /* TG68KdotC_Kernel.vhd:788:63  */
  assign n622 = n618 | n621;
  /* TG68KdotC_Kernel.vhd:788:33  */
  assign n623 = n622 ? last_data_read : ea_data;
  /* TG68KdotC_Kernel.vhd:786:33  */
  assign n624 = n617 ? addr : n623;
  /* TG68KdotC_Kernel.vhd:784:33  */
  assign n625 = n616 ? data_read : n624;
  /* TG68KdotC_Kernel.vhd:794:43  */
  assign n626 = exec[25]; // extract
  /* TG68KdotC_Kernel.vhd:797:50  */
  assign n628 = micro_state == 7'b0110010;
  /* TG68KdotC_Kernel.vhd:800:66  */
  assign n629 = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:800:87  */
  assign n630 = exec[43]; // extract
  /* TG68KdotC_Kernel.vhd:800:80  */
  assign n631 = n629 | n630;
  /* TG68KdotC_Kernel.vhd:800:98  */
  assign n632 = n631 | z_error;
  /* TG68KdotC_Kernel.vhd:801:51  */
  assign n634 = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:807:100  */
  assign n635 = trap_vector[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:807:87  */
  assign n637 = {4'b0010, n635};
  /* TG68KdotC_Kernel.vhd:809:100  */
  assign n638 = trap_vector[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:809:87  */
  assign n640 = {4'b0000, n638};
  /* TG68KdotC_Kernel.vhd:810:74  */
  assign n641 = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:810:95  */
  assign n642 = exec[43]; // extract
  /* TG68KdotC_Kernel.vhd:810:88  */
  assign n643 = n641 | n642;
  /* TG68KdotC_Kernel.vhd:810:106  */
  assign n644 = n643 | z_error;
  /* TG68KdotC_Kernel.vhd:805:41  */
  assign n645 = usestackframe2 ? n637 : n640;
  /* TG68KdotC_Kernel.vhd:805:41  */
  assign n646 = usestackframe2 ? n608 : n644;
  /* TG68KdotC_Kernel.vhd:815:43  */
  assign n647 = exec[64]; // extract
  /* TG68KdotC_Kernel.vhd:817:43  */
  assign n648 = exec[61]; // extract
  /* TG68KdotC_Kernel.vhd:819:43  */
  assign n649 = exec[62]; // extract
  /* TG68KdotC_Kernel.vhd:819:60  */
  assign n650 = ea_only & n649;
  /* TG68KdotC_Kernel.vhd:823:65  */
  assign n652 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:823:56  */
  assign n653 = n652 & exec_direct;
  /* TG68KdotC_Kernel.vhd:825:49  */
  assign n654 = exec[37]; // extract
  /* TG68KdotC_Kernel.vhd:826:94  */
  assign n655 = data_write_tmp[23:0]; // extract
  assign n656 = data_read[31:8]; // extract
  /* TG68KdotC_Kernel.vhd:825:41  */
  assign n657 = n654 ? n655 : n656;
  assign n658 = data_read[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:828:43  */
  assign n659 = exec[37]; // extract
  /* TG68KdotC_Kernel.vhd:829:78  */
  assign n660 = reg_qb[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:833:91  */
  assign n661 = {trap_sr, flags};
  assign n662 = op2out[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:832:33  */
  assign n663 = writesr ? n661 : n662;
  assign n664 = op2out[31:16]; // extract
  assign n665 = data_write_tmp[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:832:33  */
  assign n666 = writesr ? n665 : n664;
  assign n667 = {n666, n663};
  /* TG68KdotC_Kernel.vhd:830:33  */
  assign n668 = direct_data ? last_data_read : n667;
  assign n669 = n668[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:828:33  */
  assign n670 = n659 ? n660 : n669;
  assign n671 = n668[31:16]; // extract
  assign n672 = data_write_tmp[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:828:33  */
  assign n673 = n659 ? n672 : n671;
  assign n674 = {n673, n670};
  assign n675 = {n657, n658};
  /* TG68KdotC_Kernel.vhd:823:33  */
  assign n676 = n653 ? n675 : n674;
  /* TG68KdotC_Kernel.vhd:821:33  */
  assign n677 = execopc ? aluout : n676;
  /* TG68KdotC_Kernel.vhd:819:33  */
  assign n678 = n650 ? addr : n677;
  /* TG68KdotC_Kernel.vhd:817:33  */
  assign n679 = n648 ? op1out : n678;
  /* TG68KdotC_Kernel.vhd:815:33  */
  assign n680 = n647 ? data_write_tmp : n679;
  assign n681 = n680[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:801:33  */
  assign n682 = n634 ? n645 : n681;
  assign n683 = n680[31:16]; // extract
  assign n684 = data_write_tmp[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:801:33  */
  assign n685 = n634 ? n684 : n683;
  /* TG68KdotC_Kernel.vhd:801:33  */
  assign n686 = n634 ? n646 : n608;
  assign n687 = {n685, n682};
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n688 = n628 ? exe_pc : n687;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n689 = n628 ? n632 : n686;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n692 = n628 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n693 = n626 ? tg68_pc_add : n688;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n694 = n626 ? n608 : n689;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n696 = n626 ? 1'b0 : n692;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n697 = writepc ? tg68_pc : n693;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n698 = writepc ? n608 : n694;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n700 = writepc ? 1'b0 : n696;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n702 = clkena_lw ? n625 : ea_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n703 = clkena_lw ? n697 : data_write_tmp;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n704 = clkena_lw ? n606 : store_in_tmp;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n705 = clkena_lw ? n698 : writepcnext;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n706 = clkena_lw ? n585 : exec_direct;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n707 = clkena_lw ? n609 : use_direct_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n708 = clkena_lw ? n583 : direct_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n709 = clkena_lw ? n700 : usestackframe2;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n710 = clkena_lw ? n611 : z_error;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n711 = reset ? ea_data : n702;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n712 = reset ? data_write_tmp : n703;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n714 = reset ? 1'b0 : n704;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n716 = reset ? 1'b0 : n705;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n717 = reset ? exec_direct : n706;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n719 = reset ? 1'b0 : n707;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n721 = reset ? 1'b0 : n708;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n722 = reset ? usestackframe2 : n709;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n724 = reset ? 1'b0 : n710;
  /* TG68KdotC_Kernel.vhd:846:25  */
  assign n737 = brief[11]; // extract
  /* TG68KdotC_Kernel.vhd:847:46  */
  assign n738 = op1out[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n739 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n740 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n741 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n742 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n743 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n744 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n745 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n746 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n747 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n748 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n749 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n750 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n751 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n752 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n753 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:849:55  */
  assign n754 = op1out[15]; // extract
  assign n755 = {n739, n740, n741, n742};
  assign n756 = {n743, n744, n745, n746};
  assign n757 = {n747, n748, n749, n750};
  assign n758 = {n751, n752, n753, n754};
  assign n759 = {n755, n756, n757, n758};
  /* TG68KdotC_Kernel.vhd:846:17  */
  assign n760 = n737 ? n738 : n759;
  /* TG68KdotC_Kernel.vhd:851:48  */
  assign n761 = op1out[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:851:41  */
  assign n762 = {op1outbrief, n761};
  /* TG68KdotC_Kernel.vhd:852:42  */
  assign n763 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:852:50  */
  assign n765 = 1'b1 & n763;
  /* TG68KdotC_Kernel.vhd:852:35  */
  assign n767 = 1'b0 | n765;
  /* TG68KdotC_Kernel.vhd:853:35  */
  assign n768 = brief[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:854:77  */
  assign n769 = op1out[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:854:70  */
  assign n770 = {op1outbrief, n769};
  /* TG68KdotC_Kernel.vhd:854:33  */
  assign n772 = n768 == 2'b00;
  /* TG68KdotC_Kernel.vhd:855:70  */
  assign n773 = op1outbrief[14:0]; // extract
  /* TG68KdotC_Kernel.vhd:855:90  */
  assign n774 = op1out[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:855:83  */
  assign n775 = {n773, n774};
  /* TG68KdotC_Kernel.vhd:855:103  */
  assign n777 = {n775, 1'b0};
  /* TG68KdotC_Kernel.vhd:855:33  */
  assign n779 = n768 == 2'b01;
  /* TG68KdotC_Kernel.vhd:856:70  */
  assign n780 = op1outbrief[13:0]; // extract
  /* TG68KdotC_Kernel.vhd:856:90  */
  assign n781 = op1out[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:856:83  */
  assign n782 = {n780, n781};
  /* TG68KdotC_Kernel.vhd:856:103  */
  assign n784 = {n782, 2'b00};
  /* TG68KdotC_Kernel.vhd:856:33  */
  assign n786 = n768 == 2'b10;
  /* TG68KdotC_Kernel.vhd:857:70  */
  assign n787 = op1outbrief[12:0]; // extract
  /* TG68KdotC_Kernel.vhd:857:90  */
  assign n788 = op1out[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:857:83  */
  assign n789 = {n787, n788};
  /* TG68KdotC_Kernel.vhd:857:103  */
  assign n791 = {n789, 3'b000};
  /* TG68KdotC_Kernel.vhd:857:33  */
  assign n793 = n768 == 2'b11;
  assign n794 = {n793, n786, n779, n772};
  /* TG68KdotC_Kernel.vhd:853:25  */
  always @*
    case (n794)
      4'b1000: n795 = n791;
      4'b0100: n795 = n784;
      4'b0010: n795 = n777;
      4'b0001: n795 = n770;
      default: n795 = n762;
    endcase
  /* TG68KdotC_Kernel.vhd:852:17  */
  assign n796 = n767 ? n795 : n762;
  assign n803 = trap_vector[9:0]; // extract
  /* TG68KdotC_Kernel.vhd:873:33  */
  assign n804 = trap_berr ? 10'b0000001000 : n803;
  /* TG68KdotC_Kernel.vhd:876:33  */
  assign n806 = trap_addr_error ? 10'b0000001100 : n804;
  /* TG68KdotC_Kernel.vhd:879:33  */
  assign n808 = trap_illegal ? 10'b0000010000 : n806;
  /* TG68KdotC_Kernel.vhd:882:33  */
  assign n810 = set_z_error ? 10'b0000010100 : n808;
  /* TG68KdotC_Kernel.vhd:885:40  */
  assign n811 = exec[43]; // extract
  /* TG68KdotC_Kernel.vhd:885:33  */
  assign n813 = n811 ? 10'b0000011000 : n810;
  /* TG68KdotC_Kernel.vhd:888:33  */
  assign n815 = trap_trapv ? 10'b0000011100 : n813;
  /* TG68KdotC_Kernel.vhd:891:33  */
  assign n817 = trap_priv ? 10'b0000100000 : n815;
  /* TG68KdotC_Kernel.vhd:894:33  */
  assign n819 = trap_trace ? 10'b0000100100 : n817;
  /* TG68KdotC_Kernel.vhd:897:33  */
  assign n821 = trap_1010 ? 10'b0000101000 : n819;
  /* TG68KdotC_Kernel.vhd:900:33  */
  assign n823 = trap_1111 ? 10'b0000101100 : n821;
  /* TG68KdotC_Kernel.vhd:904:83  */
  assign n824 = opcode[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:904:75  */
  assign n826 = {4'b0010, n824};
  /* TG68KdotC_Kernel.vhd:904:96  */
  assign n828 = {n826, 2'b00};
  /* TG68KdotC_Kernel.vhd:903:33  */
  assign n829 = trap_trap ? n828 : n823;
  /* TG68KdotC_Kernel.vhd:906:55  */
  assign n830 = trap_interrupt | set_vectoraddr;
  /* TG68KdotC_Kernel.vhd:907:76  */
  assign n832 = {ipl_vec, 2'b00};
  /* TG68KdotC_Kernel.vhd:906:33  */
  assign n833 = n830 ? n832 : n829;
  assign n834 = {22'b0000000000000000000000, n833};
  /* TG68KdotC_Kernel.vhd:912:55  */
  assign n837 = trap_vector + vbr;
  /* TG68KdotC_Kernel.vhd:911:17  */
  assign n838 = use_vbr_stackframe ? n837 : trap_vector;
  /* TG68KdotC_Kernel.vhd:918:60  */
  assign n840 = memaddr_a[4]; // extract
  /* TG68KdotC_Kernel.vhd:918:60  */
  assign n841 = memaddr_a[4]; // extract
  /* TG68KdotC_Kernel.vhd:918:60  */
  assign n842 = memaddr_a[4]; // extract
  assign n843 = {n840, n841, n842};
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n844 = memaddr_a[7]; // extract
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n845 = memaddr_a[7]; // extract
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n846 = memaddr_a[7]; // extract
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n847 = memaddr_a[7]; // extract
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n848 = memaddr_a[7]; // extract
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n849 = memaddr_a[7]; // extract
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n850 = memaddr_a[7]; // extract
  /* TG68KdotC_Kernel.vhd:919:61  */
  assign n851 = memaddr_a[7]; // extract
  assign n852 = {n844, n845, n846, n847};
  assign n853 = {n848, n849, n850, n851};
  assign n854 = {n852, n853};
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n855 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n856 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n857 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n858 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n859 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n860 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n861 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n862 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n863 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n864 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n865 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n866 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n867 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n868 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n869 = memaddr_a[15]; // extract
  /* TG68KdotC_Kernel.vhd:920:62  */
  assign n870 = memaddr_a[15]; // extract
  assign n871 = {n855, n856, n857, n858};
  assign n872 = {n859, n860, n861, n862};
  assign n873 = {n863, n864, n865, n866};
  assign n874 = {n867, n868, n869, n870};
  assign n875 = {n871, n872, n873, n874};
  /* TG68KdotC_Kernel.vhd:922:32  */
  assign n876 = exec[70]; // extract
  /* TG68KdotC_Kernel.vhd:923:55  */
  assign n877 = briefdata + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:925:72  */
  assign n878 = last_data_read[7:0]; // extract
  assign n879 = last_data_read[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:924:25  */
  assign n880 = setdispbyte ? n878 : n879;
  assign n881 = last_data_read[31:8]; // extract
  assign n882 = {n875, n854};
  /* TG68KdotC_Kernel.vhd:924:25  */
  assign n883 = setdispbyte ? n882 : n881;
  assign n884 = {n883, n880};
  /* TG68KdotC_Kernel.vhd:922:25  */
  assign n885 = n876 ? n877 : n884;
  /* TG68KdotC_Kernel.vhd:929:26  */
  assign n886 = set[47]; // extract
  /* TG68KdotC_Kernel.vhd:930:31  */
  assign n887 = set[73]; // extract
  /* TG68KdotC_Kernel.vhd:932:39  */
  assign n890 = datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:932:52  */
  assign n891 = set[50]; // extract
  /* TG68KdotC_Kernel.vhd:932:60  */
  assign n892 = ~n891;
  /* TG68KdotC_Kernel.vhd:932:45  */
  assign n893 = n892 & n890;
  /* TG68KdotC_Kernel.vhd:932:25  */
  assign n896 = n893 ? 5'b11111 : 5'b11110;
  /* TG68KdotC_Kernel.vhd:930:25  */
  assign n897 = n887 ? 5'b11100 : n896;
  /* TG68KdotC_Kernel.vhd:938:53  */
  assign n899 = {1'b1, ripl_nr};
  /* TG68KdotC_Kernel.vhd:938:61  */
  assign n901 = {n899, 1'b0};
  /* TG68KdotC_Kernel.vhd:937:17  */
  assign n902 = interrupt ? n901 : 5'b00000;
  /* TG68KdotC_Kernel.vhd:929:17  */
  assign n903 = n886 ? n897 : n902;
  assign n904 = n885[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:921:17  */
  assign n905 = setdisp ? n904 : n903;
  assign n906 = n885[31:5]; // extract
  assign n907 = {n875, n854, n843};
  /* TG68KdotC_Kernel.vhd:921:17  */
  assign n908 = setdisp ? n906 : n907;
  /* TG68KdotC_Kernel.vhd:943:40  */
  assign n910 = exec[71]; // extract
  /* TG68KdotC_Kernel.vhd:943:66  */
  assign n912 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:943:83  */
  assign n913 = memread[0]; // extract
  /* TG68KdotC_Kernel.vhd:943:72  */
  assign n914 = n913 & n912;
  /* TG68KdotC_Kernel.vhd:943:57  */
  assign n915 = n910 | n914;
  /* TG68KdotC_Kernel.vhd:948:46  */
  assign n917 = memmaskmux[3]; // extract
  /* TG68KdotC_Kernel.vhd:948:49  */
  assign n918 = ~n917;
  /* TG68KdotC_Kernel.vhd:948:61  */
  assign n919 = exec[55]; // extract
  /* TG68KdotC_Kernel.vhd:948:54  */
  assign n920 = n918 | n919;
  /* TG68KdotC_Kernel.vhd:950:42  */
  assign n921 = set[83]; // extract
  /* TG68KdotC_Kernel.vhd:952:43  */
  assign n922 = exec[58]; // extract
  /* TG68KdotC_Kernel.vhd:954:43  */
  assign n923 = exec[63]; // extract
  /* TG68KdotC_Kernel.vhd:954:70  */
  assign n925 = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:954:58  */
  assign n926 = n925 & n923;
  /* TG68KdotC_Kernel.vhd:956:42  */
  assign n927 = set[45]; // extract
  /* TG68KdotC_Kernel.vhd:958:47  */
  assign n929 = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:960:43  */
  assign n930 = exec[22]; // extract
  /* TG68KdotC_Kernel.vhd:967:53  */
  assign n931 = ~interrupt;
  /* TG68KdotC_Kernel.vhd:967:75  */
  assign n932 = ~suppress_base;
  /* TG68KdotC_Kernel.vhd:967:58  */
  assign n933 = n932 & n931;
  /* TG68KdotC_Kernel.vhd:967:41  */
  assign n936 = n933 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:963:33  */
  assign n937 = set_vectoraddr ? trap_vector_vbr : memaddr_a;
  /* TG68KdotC_Kernel.vhd:963:33  */
  assign n939 = set_vectoraddr ? 1'b0 : n936;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n940 = n930 ? ea_data : n937;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n942 = n930 ? memaddr_a : 32'b00000000000000000000000000000000;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n944 = n930 ? 1'b0 : n939;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n945 = n929 ? tg68_pc_add : n940;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n947 = n929 ? 32'b00000000000000000000000000000000 : n942;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n949 = n929 ? 1'b0 : n944;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n950 = n927 ? last_data_read : n945;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n952 = n927 ? 32'b00000000000000000000000000000000 : n947;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n954 = n927 ? 1'b0 : n949;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n955 = n926 ? addr : n950;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n957 = n926 ? 32'b00000000000000000000000000000000 : n952;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n959 = n926 ? 1'b0 : n954;
  /* TG68KdotC_Kernel.vhd:952:33  */
  assign n960 = n922 ? data_read : n955;
  /* TG68KdotC_Kernel.vhd:952:33  */
  assign n962 = n922 ? 32'b00000000000000000000000000000000 : n957;
  /* TG68KdotC_Kernel.vhd:952:33  */
  assign n964 = n922 ? 1'b0 : n959;
  /* TG68KdotC_Kernel.vhd:950:33  */
  assign n965 = n921 ? tmp_tg68_pc : n960;
  /* TG68KdotC_Kernel.vhd:950:33  */
  assign n967 = n921 ? 32'b00000000000000000000000000000000 : n962;
  /* TG68KdotC_Kernel.vhd:950:33  */
  assign n969 = n921 ? 1'b0 : n964;
  /* TG68KdotC_Kernel.vhd:948:33  */
  assign n970 = n920 ? addsub_q : n965;
  /* TG68KdotC_Kernel.vhd:948:33  */
  assign n972 = n920 ? 32'b00000000000000000000000000000000 : n967;
  /* TG68KdotC_Kernel.vhd:948:33  */
  assign n975 = n920 ? 1'b0 : n969;
  /* TG68KdotC_Kernel.vhd:975:53  */
  assign n977 = memread[0]; // extract
  /* TG68KdotC_Kernel.vhd:975:73  */
  assign n978 = state[1]; // extract
  /* TG68KdotC_Kernel.vhd:975:64  */
  assign n979 = n978 & n977;
  /* TG68KdotC_Kernel.vhd:975:100  */
  assign n980 = ~movem_presub;
  /* TG68KdotC_Kernel.vhd:975:84  */
  assign n981 = n979 | n980;
  /* TG68KdotC_Kernel.vhd:942:25  */
  assign n983 = n915 & clkena_in;
  /* TG68KdotC_Kernel.vhd:942:25  */
  assign n984 = n981 & clkena_in;
  /* TG68KdotC_Kernel.vhd:981:53  */
  assign n993 = memaddr_delta_rega + memaddr_delta_regb;
  /* TG68KdotC_Kernel.vhd:983:36  */
  assign n994 = memaddr_reg + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:984:41  */
  assign n995 = memaddr_reg + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:986:28  */
  assign n996 = ~use_base;
  /* TG68KdotC_Kernel.vhd:986:17  */
  assign n998 = n996 ? 32'b00000000000000000000000000000000 : reg_qa;
  /* TG68KdotC_Kernel.vhd:1001:17  */
  assign n1002 = tg68_pc_brw ? tmp_tg68_pc : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1006:40  */
  assign n1004 = pc_datab[2]; // extract
  /* TG68KdotC_Kernel.vhd:1007:60  */
  assign n1005 = pc_datab[3]; // extract
  /* TG68KdotC_Kernel.vhd:1007:60  */
  assign n1006 = pc_datab[3]; // extract
  /* TG68KdotC_Kernel.vhd:1007:60  */
  assign n1007 = pc_datab[3]; // extract
  /* TG68KdotC_Kernel.vhd:1007:60  */
  assign n1008 = pc_datab[3]; // extract
  assign n1009 = {n1005, n1006, n1007, n1008};
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1010 = pc_datab[7]; // extract
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1011 = pc_datab[7]; // extract
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1012 = pc_datab[7]; // extract
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1013 = pc_datab[7]; // extract
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1014 = pc_datab[7]; // extract
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1015 = pc_datab[7]; // extract
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1016 = pc_datab[7]; // extract
  /* TG68KdotC_Kernel.vhd:1008:61  */
  assign n1017 = pc_datab[7]; // extract
  assign n1018 = {n1010, n1011, n1012, n1013};
  assign n1019 = {n1014, n1015, n1016, n1017};
  assign n1020 = {n1018, n1019};
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1021 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1022 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1023 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1024 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1025 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1026 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1027 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1028 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1029 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1030 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1031 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1032 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1033 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1034 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1035 = pc_datab[15]; // extract
  /* TG68KdotC_Kernel.vhd:1009:62  */
  assign n1036 = pc_datab[15]; // extract
  assign n1037 = {n1021, n1022, n1023, n1024};
  assign n1038 = {n1025, n1026, n1027, n1028};
  assign n1039 = {n1029, n1030, n1031, n1032};
  assign n1040 = {n1033, n1034, n1035, n1036};
  assign n1041 = {n1037, n1038, n1039, n1040};
  assign n1043 = n1003[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1010:17  */
  assign n1044 = interrupt ? 2'b11 : n1043;
  assign n1045 = n1003[0]; // extract
  /* TG68KdotC_Kernel.vhd:1013:24  */
  assign n1046 = exec[25]; // extract
  assign n1050 = n1044[0]; // extract
  /* TG68KdotC_Kernel.vhd:1014:25  */
  assign n1051 = writepcbig ? 1'b1 : n1050;
  assign n1052 = n1044[1]; // extract
  /* TG68KdotC_Kernel.vhd:1014:25  */
  assign n1053 = writepcbig ? n1052 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1014:25  */
  assign n1054 = writepcbig ? 1'b1 : n1004;
  /* TG68KdotC_Kernel.vhd:1020:47  */
  assign n1055 = ~use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:1020:71  */
  assign n1056 = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:1020:96  */
  assign n1057 = exec[43]; // extract
  /* TG68KdotC_Kernel.vhd:1020:89  */
  assign n1058 = n1056 | n1057;
  /* TG68KdotC_Kernel.vhd:1020:111  */
  assign n1059 = n1058 | z_error;
  /* TG68KdotC_Kernel.vhd:1020:52  */
  assign n1060 = n1059 & n1055;
  /* TG68KdotC_Kernel.vhd:1020:128  */
  assign n1061 = n1060 | writepcnext;
  /* TG68KdotC_Kernel.vhd:1020:25  */
  assign n1063 = n1061 ? 1'b1 : n1051;
  /* TG68KdotC_Kernel.vhd:1023:28  */
  assign n1065 = state == 2'b00;
  assign n1067 = n1044[0]; // extract
  /* TG68KdotC_Kernel.vhd:1023:17  */
  assign n1068 = n1065 ? 1'b1 : n1067;
  assign n1069 = {n1054, n1053, n1063};
  assign n1070 = n1069[0]; // extract
  /* TG68KdotC_Kernel.vhd:1013:17  */
  assign n1071 = n1046 ? n1070 : n1068;
  assign n1072 = n1069[2:1]; // extract
  assign n1073 = n1044[1]; // extract
  assign n1074 = {n1004, n1073};
  /* TG68KdotC_Kernel.vhd:1013:17  */
  assign n1075 = n1046 ? n1072 : n1074;
  /* TG68KdotC_Kernel.vhd:1030:63  */
  assign n1077 = opcode[7:0]; // extract
  assign n1078 = last_data_read[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:1027:25  */
  assign n1079 = tg68_pc_word ? n1078 : n1077;
  assign n1080 = last_data_read[31:8]; // extract
  assign n1081 = {n1041, n1020};
  /* TG68KdotC_Kernel.vhd:1027:25  */
  assign n1082 = tg68_pc_word ? n1080 : n1081;
  assign n1083 = {n1082, n1079};
  assign n1084 = {n1041, n1020, n1009, n1075, n1071, n1045};
  /* TG68KdotC_Kernel.vhd:1026:17  */
  assign n1085 = tg68_pc_brw ? n1083 : n1084;
  /* TG68KdotC_Kernel.vhd:1034:40  */
  assign n1086 = pc_dataa + pc_datab;
  /* TG68KdotC_Kernel.vhd:1039:28  */
  assign n1088 = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1039:54  */
  assign n1090 = next_micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1039:34  */
  assign n1091 = n1090 & n1088;
  /* TG68KdotC_Kernel.vhd:1039:75  */
  assign n1092 = ~setnextpass;
  /* TG68KdotC_Kernel.vhd:1039:60  */
  assign n1093 = n1092 & n1091;
  /* TG68KdotC_Kernel.vhd:1039:100  */
  assign n1094 = ~exec_write_back;
  /* TG68KdotC_Kernel.vhd:1039:113  */
  assign n1096 = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:1039:105  */
  assign n1097 = n1094 | n1096;
  /* TG68KdotC_Kernel.vhd:1039:80  */
  assign n1098 = n1097 & n1093;
  /* TG68KdotC_Kernel.vhd:1039:135  */
  assign n1100 = set_rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:1039:120  */
  assign n1101 = n1100 & n1098;
  /* TG68KdotC_Kernel.vhd:1039:157  */
  assign n1102 = set_exec[31]; // extract
  /* TG68KdotC_Kernel.vhd:1039:165  */
  assign n1103 = ~n1102;
  /* TG68KdotC_Kernel.vhd:1039:145  */
  assign n1104 = n1103 & n1101;
  /* TG68KdotC_Kernel.vhd:1041:35  */
  assign n1105 = flagssr[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1041:47  */
  assign n1106 = $unsigned(n1105) < $unsigned(ipl_nr);
  /* TG68KdotC_Kernel.vhd:1041:64  */
  assign n1108 = ipl_nr == 3'b111;
  /* TG68KdotC_Kernel.vhd:1041:55  */
  assign n1109 = n1106 | n1108;
  /* TG68KdotC_Kernel.vhd:1041:72  */
  assign n1110 = n1109 | make_trace;
  /* TG68KdotC_Kernel.vhd:1041:90  */
  assign n1111 = n1110 | make_berr;
  /* TG68KdotC_Kernel.vhd:1043:35  */
  assign n1112 = ~stop;
  /* TG68KdotC_Kernel.vhd:1043:25  */
  assign n1115 = n1112 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1041:25  */
  assign n1117 = n1111 ? 1'b0 : n1115;
  /* TG68KdotC_Kernel.vhd:1041:25  */
  assign n1120 = n1111 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1039:17  */
  assign n1122 = n1104 ? n1117 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1039:17  */
  assign n1126 = n1104 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1039:17  */
  assign n1129 = n1104 ? n1120 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1048:28  */
  assign n1132 = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1048:54  */
  assign n1134 = next_micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1048:34  */
  assign n1135 = n1134 & n1132;
  /* TG68KdotC_Kernel.vhd:1048:79  */
  assign n1136 = ~set_direct_data;
  /* TG68KdotC_Kernel.vhd:1048:60  */
  assign n1137 = n1136 & n1135;
  /* TG68KdotC_Kernel.vhd:1048:104  */
  assign n1138 = ~exec_write_back;
  /* TG68KdotC_Kernel.vhd:1048:118  */
  assign n1140 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1048:137  */
  assign n1141 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:1048:124  */
  assign n1142 = n1141 & n1140;
  /* TG68KdotC_Kernel.vhd:1048:109  */
  assign n1143 = n1138 | n1142;
  /* TG68KdotC_Kernel.vhd:1048:84  */
  assign n1144 = n1143 & n1137;
  /* TG68KdotC_Kernel.vhd:1048:17  */
  assign n1147 = n1144 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1052:27  */
  assign n1149 = ~IPL;
  /* TG68KdotC_Kernel.vhd:1082:59  */
  assign n1151 = memmask[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:1082:71  */
  assign n1153 = {n1151, 2'b11};
  /* TG68KdotC_Kernel.vhd:1083:59  */
  assign n1154 = memread[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:1083:82  */
  assign n1155 = memmaskmux[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1083:71  */
  assign n1156 = {n1154, n1155};
  /* TG68KdotC_Kernel.vhd:1087:48  */
  assign n1157 = exec[57]; // extract
  /* TG68KdotC_Kernel.vhd:1089:51  */
  assign n1158 = exec[63]; // extract
  /* TG68KdotC_Kernel.vhd:1091:54  */
  assign n1160 = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1091:60  */
  assign n1161 = n1160 | tg68_pc_brw;
  /* TG68KdotC_Kernel.vhd:1091:90  */
  assign n1162 = ~stop;
  /* TG68KdotC_Kernel.vhd:1091:82  */
  assign n1163 = n1162 & n1161;
  /* TG68KdotC_Kernel.vhd:1091:41  */
  assign n1164 = n1163 ? tg68_pc_add : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1089:41  */
  assign n1165 = n1158 ? addr : n1164;
  /* TG68KdotC_Kernel.vhd:1087:41  */
  assign n1166 = n1157 ? data_read : n1165;
  /* TG68KdotC_Kernel.vhd:1081:33  */
  assign n1167 = clkena_in ? n1166 : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1081:33  */
  assign n1168 = clkena_in ? n1153 : memmask;
  /* TG68KdotC_Kernel.vhd:1081:33  */
  assign n1169 = clkena_in ? n1156 : memread;
  /* TG68KdotC_Kernel.vhd:1109:53  */
  assign n1170 = ~trap_berr;
  /* TG68KdotC_Kernel.vhd:1110:68  */
  assign n1171 = berr | make_berr;
  /* TG68KdotC_Kernel.vhd:1109:41  */
  assign n1173 = n1170 ? n1171 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1115:71  */
  assign n1174 = ~setinterrupt;
  /* TG68KdotC_Kernel.vhd:1115:67  */
  assign n1175 = n1174 & stop;
  /* TG68KdotC_Kernel.vhd:1115:58  */
  assign n1176 = set_stop | n1175;
  /* TG68KdotC_Kernel.vhd:1128:75  */
  assign n1178 = {5'b00011, ipl_nr};
  /* TG68KdotC_Kernel.vhd:1124:49  */
  assign n1181 = make_berr ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1124:49  */
  assign n1184 = make_berr ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1124:49  */
  assign n1185 = make_berr ? ripl_nr : ipl_nr;
  /* TG68KdotC_Kernel.vhd:1124:49  */
  assign n1186 = make_berr ? ipl_vec : n1178;
  /* TG68KdotC_Kernel.vhd:1122:49  */
  assign n1188 = make_trace ? 1'b0 : n1181;
  /* TG68KdotC_Kernel.vhd:1122:49  */
  assign n1192 = make_trace ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1122:49  */
  assign n1195 = make_trace ? 1'b0 : n1184;
  /* TG68KdotC_Kernel.vhd:1122:49  */
  assign n1197 = make_trace ? ripl_nr : n1185;
  /* TG68KdotC_Kernel.vhd:1122:49  */
  assign n1198 = make_trace ? ipl_vec : n1186;
  /* TG68KdotC_Kernel.vhd:1116:41  */
  assign n1199 = setinterrupt ? n1188 : trap_berr;
  /* TG68KdotC_Kernel.vhd:1116:41  */
  assign n1200 = setinterrupt ? n1192 : trap_trace;
  /* TG68KdotC_Kernel.vhd:1116:41  */
  assign n1201 = setinterrupt ? n1195 : trap_interrupt;
  /* TG68KdotC_Kernel.vhd:1116:41  */
  assign n1203 = setinterrupt ? 1'b0 : n1173;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1204 = n1407 ? n1197 : ripl_nr;
  /* TG68KdotC_Kernel.vhd:1116:41  */
  assign n1205 = setinterrupt ? n1198 : ipl_vec;
  /* TG68KdotC_Kernel.vhd:1132:55  */
  assign n1207 = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1132:80  */
  assign n1208 = ~IPL_autovector;
  /* TG68KdotC_Kernel.vhd:1132:62  */
  assign n1209 = n1208 & n1207;
  /* TG68KdotC_Kernel.vhd:1133:74  */
  assign n1210 = last_data_read[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:1132:41  */
  assign n1211 = n1209 ? n1210 : n1205;
  /* TG68KdotC_Kernel.vhd:1135:49  */
  assign n1213 = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1136:75  */
  assign n1214 = data_read[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1215 = n1389 ? tg68_pc : last_opc_pc;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1216 = n1390 ? n1214 : last_opc_read;
  /* TG68KdotC_Kernel.vhd:1144:53  */
  assign n1217 = opcode[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:1144:65  */
  assign n1219 = n1217 == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:1144:86  */
  assign n1220 = opcode[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:1144:98  */
  assign n1222 = n1220 == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:1144:77  */
  assign n1223 = n1219 | n1222;
  /* TG68KdotC_Kernel.vhd:1144:110  */
  assign n1224 = n1223 | data_is_source;
  /* TG68KdotC_Kernel.vhd:1144:41  */
  assign n1226 = n1224 ? 1'b1 : tg68_pc_word;
  /* TG68KdotC_Kernel.vhd:1139:41  */
  assign n1228 = setopcode ? 1'b0 : n1226;
  /* TG68KdotC_Kernel.vhd:1139:41  */
  assign n1230 = setopcode ? 1'b0 : n1199;
  /* TG68KdotC_Kernel.vhd:1139:41  */
  assign n1232 = setopcode ? 1'b0 : n1200;
  /* TG68KdotC_Kernel.vhd:1139:41  */
  assign n1234 = setopcode ? 1'b0 : n1201;
  /* TG68KdotC_Kernel.vhd:1148:48  */
  assign n1235 = exec[29]; // extract
  /* TG68KdotC_Kernel.vhd:1152:84  */
  assign n1236 = {26'b0, bf_width};  //  uext
  /* TG68KdotC_Kernel.vhd:1152:84  */
  assign n1237 = bf_full_offset + n1236;
  /* TG68KdotC_Kernel.vhd:1152:93  */
  assign n1239 = n1237 + 32'b00000000000000000000000000000001;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1240 = n1416 ? bf_width : alu_width;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1241 = n1417 ? bf_shift : alu_bf_shift;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1242 = n1418 ? n1239 : alu_bf_ffo_offset;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1243 = n1419 ? bf_loffset : alu_bf_loffset;
  /* TG68KdotC_Kernel.vhd:1155:62  */
  assign n1244 = setstate[1]; // extract
  /* TG68KdotC_Kernel.vhd:1155:50  */
  assign n1245 = ~n1244;
  /* TG68KdotC_Kernel.vhd:1155:93  */
  assign n1246 = setstate[0]; // extract
  /* TG68KdotC_Kernel.vhd:1155:81  */
  assign n1247 = ~n1246;
  /* TG68KdotC_Kernel.vhd:1155:77  */
  assign n1248 = pcbase & n1247;
  /* TG68KdotC_Kernel.vhd:1155:66  */
  assign n1249 = n1245 | n1248;
  /* TG68KdotC_Kernel.vhd:1156:58  */
  assign n1250 = setstate[1]; // extract
  /* TG68KdotC_Kernel.vhd:1156:67  */
  assign n1251 = ~pcbase;
  /* TG68KdotC_Kernel.vhd:1156:89  */
  assign n1252 = setstate[0]; // extract
  /* TG68KdotC_Kernel.vhd:1156:78  */
  assign n1253 = n1251 | n1252;
  /* TG68KdotC_Kernel.vhd:1156:62  */
  assign n1254 = n1250 & n1253;
  assign n1256 = {n1249, n1254};
  /* TG68KdotC_Kernel.vhd:1157:41  */
  assign n1257 = interrupt ? 2'b11 : n1256;
  /* TG68KdotC_Kernel.vhd:1161:49  */
  assign n1259 = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:1163:55  */
  assign n1261 = setstate == 2'b10;
  /* TG68KdotC_Kernel.vhd:1163:77  */
  assign n1262 = ~setaddrvalue;
  /* TG68KdotC_Kernel.vhd:1163:61  */
  assign n1263 = n1262 & n1261;
  /* TG68KdotC_Kernel.vhd:1163:82  */
  assign n1264 = write_back & n1263;
  /* TG68KdotC_Kernel.vhd:1163:41  */
  assign n1266 = n1264 ? 1'b1 : exec_write_back;
  /* TG68KdotC_Kernel.vhd:1161:41  */
  assign n1268 = n1259 ? 1'b0 : n1266;
  /* TG68KdotC_Kernel.vhd:1166:50  */
  assign n1270 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1166:69  */
  assign n1271 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:1166:56  */
  assign n1272 = n1271 & n1270;
  /* TG68KdotC_Kernel.vhd:1166:74  */
  assign n1273 = write_back & n1272;
  /* TG68KdotC_Kernel.vhd:1166:105  */
  assign n1275 = setstate != 2'b10;
  /* TG68KdotC_Kernel.vhd:1166:93  */
  assign n1276 = n1275 & n1273;
  /* TG68KdotC_Kernel.vhd:1166:127  */
  assign n1278 = set_rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1166:113  */
  assign n1279 = n1276 | n1278;
  /* TG68KdotC_Kernel.vhd:1166:164  */
  assign n1280 = ~interrupt;
  /* TG68KdotC_Kernel.vhd:1166:151  */
  assign n1281 = n1280 & stop;
  /* TG68KdotC_Kernel.vhd:1166:138  */
  assign n1282 = n1279 | n1281;
  /* TG68KdotC_Kernel.vhd:1166:181  */
  assign n1283 = set_exec[31]; // extract
  /* TG68KdotC_Kernel.vhd:1166:170  */
  assign n1284 = n1282 | n1283;
  /* TG68KdotC_Kernel.vhd:1170:59  */
  assign n1285 = exec_write_back & execopc;
  /* TG68KdotC_Kernel.vhd:1178:60  */
  assign n1288 = setstate == 2'b01;
  /* TG68KdotC_Kernel.vhd:1181:59  */
  assign n1289 = exec[29]; // extract
  /* TG68KdotC_Kernel.vhd:1185:58  */
  assign n1290 = set[73]; // extract
  /* TG68KdotC_Kernel.vhd:1190:67  */
  assign n1292 = set_datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:1190:85  */
  assign n1293 = setstate[1]; // extract
  /* TG68KdotC_Kernel.vhd:1190:73  */
  assign n1294 = n1293 & n1292;
  /* TG68KdotC_Kernel.vhd:1193:63  */
  assign n1295 = set[72]; // extract
  /* TG68KdotC_Kernel.vhd:1193:57  */
  assign n1298 = n1295 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1190:49  */
  assign n1301 = n1294 ? 6'b101111 : 6'b100111;
  /* TG68KdotC_Kernel.vhd:1190:49  */
  assign n1304 = n1294 ? 6'b101111 : 6'b100111;
  /* TG68KdotC_Kernel.vhd:1190:49  */
  assign n1306 = n1294 ? n1298 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1185:49  */
  assign n1308 = n1290 ? 6'b100001 : n1301;
  /* TG68KdotC_Kernel.vhd:1185:49  */
  assign n1310 = n1290 ? 6'b100001 : n1304;
  /* TG68KdotC_Kernel.vhd:1185:49  */
  assign n1312 = n1290 ? 1'b0 : n1306;
  /* TG68KdotC_Kernel.vhd:1181:49  */
  assign n1313 = n1289 ? set_memmask : n1308;
  /* TG68KdotC_Kernel.vhd:1181:49  */
  assign n1314 = n1289 ? set_memmask : n1310;
  /* TG68KdotC_Kernel.vhd:1181:49  */
  assign n1315 = n1289 ? set_oddout : n1312;
  /* TG68KdotC_Kernel.vhd:1178:49  */
  assign n1317 = n1288 ? 6'b111111 : n1313;
  /* TG68KdotC_Kernel.vhd:1178:49  */
  assign n1319 = n1288 ? 6'b111111 : n1314;
  /* TG68KdotC_Kernel.vhd:1178:49  */
  assign n1320 = n1288 ? oddout : n1315;
  /* TG68KdotC_Kernel.vhd:1170:41  */
  assign n1321 = n1285 ? 2'b01 : n1257;
  /* TG68KdotC_Kernel.vhd:1170:41  */
  assign n1323 = n1285 ? 2'b11 : setstate;
  /* TG68KdotC_Kernel.vhd:1170:41  */
  assign n1325 = n1285 ? 1'b0 : setaddrvalue;
  /* TG68KdotC_Kernel.vhd:1170:41  */
  assign n1326 = n1285 ? wbmemmask : n1317;
  /* TG68KdotC_Kernel.vhd:1170:41  */
  assign n1327 = n1285 ? wbmemmask : n1319;
  /* TG68KdotC_Kernel.vhd:1170:41  */
  assign n1328 = n1285 ? oddout : n1320;
  /* TG68KdotC_Kernel.vhd:1166:41  */
  assign n1329 = n1284 ? n1257 : n1321;
  /* TG68KdotC_Kernel.vhd:1166:41  */
  assign n1331 = n1284 ? 2'b01 : n1323;
  /* TG68KdotC_Kernel.vhd:1166:41  */
  assign n1333 = n1284 ? 1'b0 : n1325;
  /* TG68KdotC_Kernel.vhd:1166:41  */
  assign n1335 = n1284 ? 6'b111111 : n1326;
  /* TG68KdotC_Kernel.vhd:1166:41  */
  assign n1336 = n1284 ? wbmemmask : n1327;
  /* TG68KdotC_Kernel.vhd:1166:41  */
  assign n1337 = n1284 ? oddout : n1328;
  /* TG68KdotC_Kernel.vhd:1209:78  */
  assign n1338 = set_writepcbig | writepcbig;
  /* TG68KdotC_Kernel.vhd:1205:41  */
  assign n1340 = decodeopc ? 1'b0 : n1338;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1341 = n1399 ? set_rot_bits : rot_bits;
  /* TG68KdotC_Kernel.vhd:1211:65  */
  assign n1342 = exec[24]; // extract
  /* TG68KdotC_Kernel.vhd:1211:58  */
  assign n1343 = decodeopc | n1342;
  /* TG68KdotC_Kernel.vhd:1211:92  */
  assign n1345 = rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1211:82  */
  assign n1346 = n1343 | n1345;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1347 = n1400 ? set_rot_cnt : rot_cnt;
  /* TG68KdotC_Kernel.vhd:1217:55  */
  assign n1348 = setstate[1]; // extract
  /* TG68KdotC_Kernel.vhd:1217:86  */
  assign n1349 = set[62]; // extract
  /* TG68KdotC_Kernel.vhd:1217:79  */
  assign n1350 = n1349 & ea_only;
  /* TG68KdotC_Kernel.vhd:1217:63  */
  assign n1351 = n1348 | n1350;
  /* TG68KdotC_Kernel.vhd:1217:41  */
  assign n1353 = n1351 ? 1'b0 : suppress_base;
  /* TG68KdotC_Kernel.vhd:1215:41  */
  assign n1355 = set_suppress_base ? 1'b1 : n1353;
  /* TG68KdotC_Kernel.vhd:1221:57  */
  assign n1356 = state[1]; // extract
  /* TG68KdotC_Kernel.vhd:1224:75  */
  assign n1357 = data_read[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:1221:49  */
  assign n1358 = n1356 ? last_opc_read : n1357;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1359 = n1393 ? n1358 : brief;
  /* TG68KdotC_Kernel.vhd:1228:66  */
  assign n1360 = ~berr;
  /* TG68KdotC_Kernel.vhd:1228:58  */
  assign n1361 = n1360 & setopcode;
  /* TG68KdotC_Kernel.vhd:1229:57  */
  assign n1363 = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1230:76  */
  assign n1364 = data_read[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:1229:49  */
  assign n1365 = n1363 ? n1364 : last_opc_read;
  /* TG68KdotC_Kernel.vhd:1229:49  */
  assign n1366 = n1363 ? tg68_pc : last_opc_pc;
  /* TG68KdotC_Kernel.vhd:1237:64  */
  assign n1367 = setinterrupt | setopcode;
  /* TG68KdotC_Kernel.vhd:1242:68  */
  assign n1368 = setnextpass | regdirectsource;
  /* TG68KdotC_Kernel.vhd:1242:49  */
  assign n1370 = n1368 ? 1'b1 : nextpass;
  /* TG68KdotC_Kernel.vhd:1237:41  */
  assign n1372 = n1367 ? 16'b0100111001110001 : opcode;
  /* TG68KdotC_Kernel.vhd:1237:41  */
  assign n1374 = n1367 ? 1'b0 : n1370;
  /* TG68KdotC_Kernel.vhd:1228:41  */
  assign n1375 = n1361 ? n1365 : n1372;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1376 = n1388 ? n1366 : exe_pc;
  /* TG68KdotC_Kernel.vhd:1228:41  */
  assign n1378 = n1361 ? 1'b0 : n1374;
  /* TG68KdotC_Kernel.vhd:1247:58  */
  assign n1379 = decodeopc | interrupt;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1380 = n1404 ? flagssr : trap_sr;
  assign n1381 = n9425[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1382 = clkena_lw ? n1329 : n1381;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1383 = clkena_lw ? n1331 : state;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1384 = clkena_lw ? set_datatype : exe_datatype;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1385 = clkena_lw ? n1333 : addrvalue;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1386 = clkena_lw ? n1375 : opcode;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1387 = clkena_lw ? opcode : exe_opcode;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1388 = n1361 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1389 = n1213 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1390 = n1213 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1391 = clkena_lw ? n1378 : nextpass;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1392 = clkena_lw ? n1228 : tg68_pc_word;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1393 = getbrief & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1394 = clkena_lw ? n1268 : exec_write_back;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1395 = clkena_lw ? n1340 : writepcbig;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1396 = clkena_lw ? setopcode : decodeopc;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1397 = clkena_lw ? setexecopc : execopc;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1398 = clkena_lw ? setendopc : endopc;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1399 = decodeopc & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1400 = n1346 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1401 = clkena_lw ? n1230 : trap_berr;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1402 = clkena_lw ? n1232 : trap_trace;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1403 = clkena_lw ? n1234 : trap_interrupt;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1404 = n1379 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1405 = clkena_lw ? n1203 : make_berr;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1406 = clkena_lw ? n1176 : stop;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1407 = setinterrupt & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1408 = clkena_lw ? n1211 : ipl_vec;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1409 = clkena_lw ? setinterrupt : interrupt;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1410 = clkena_lw ? n1355 : suppress_base;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1411 = clkena_lw ? n1335 : n1168;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1413 = clkena_lw ? 4'b1111 : n1169;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1414 = clkena_lw ? n1336 : wbmemmask;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1415 = clkena_lw ? n1337 : oddout;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1416 = n1235 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1417 = n1235 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1418 = n1235 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1095:33  */
  assign n1419 = n1235 & clkena_lw;
  assign n1420 = n9425[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1421 = reset ? n1420 : n1382;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1423 = reset ? 32'b00000000000000000000000000000100 : n1167;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1425 = reset ? 2'b01 : n1383;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1426 = reset ? exe_datatype : n1384;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1428 = reset ? 1'b0 : n1385;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1430 = reset ? 16'b0010111001111001 : n1386;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1431 = reset ? exe_opcode : n1387;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1432 = reset ? exe_pc : n1376;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1433 = reset ? last_opc_pc : n1215;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1435 = reset ? 16'b0100111011111001 : n1216;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1436 = reset ? nextpass : n1391;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1438 = reset ? 1'b0 : n1392;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1439 = reset ? brief : n1359;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1441 = reset ? 1'b0 : n1394;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1443 = reset ? 1'b0 : n1395;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1445 = reset ? 1'b0 : n1396;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1447 = reset ? 1'b0 : n1397;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1449 = reset ? 1'b0 : n1398;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1450 = reset ? rot_bits : n1341;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1452 = reset ? 6'b000001 : n1347;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1454 = reset ? 1'b0 : n1401;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1456 = reset ? 1'b0 : n1402;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1458 = reset ? 1'b0 : n1403;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1459 = reset ? trap_sr : n1380;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1461 = reset ? 1'b0 : n1405;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1463 = reset ? 1'b0 : n1406;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1464 = reset ? ripl_nr : n1204;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1465 = reset ? ipl_vec : n1408;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1467 = reset ? 1'b0 : n1409;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1469 = reset ? 1'b0 : n1410;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1471 = reset ? 6'b111111 : n1411;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1472 = reset ? memread : n1413;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1473 = reset ? wbmemmask : n1414;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1474 = reset ? oddout : n1415;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1475 = reset ? alu_width : n1240;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1476 = reset ? alu_bf_shift : n1241;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1477 = reset ? alu_bf_ffo_offset : n1242;
  /* TG68KdotC_Kernel.vhd:1054:25  */
  assign n1478 = reset ? alu_bf_loffset : n1243;
  /* TG68KdotC_Kernel.vhd:1258:54  */
  assign n1519 = set_pcbase | pcbase;
  /* TG68KdotC_Kernel.vhd:1259:60  */
  assign n1520 = state[1]; // extract
  /* TG68KdotC_Kernel.vhd:1259:81  */
  assign n1521 = ~movem_run;
  /* TG68KdotC_Kernel.vhd:1259:68  */
  assign n1522 = n1521 & n1520;
  /* TG68KdotC_Kernel.vhd:1259:51  */
  assign n1523 = setexecopc | n1522;
  /* TG68KdotC_Kernel.vhd:1259:33  */
  assign n1525 = n1523 ? 1'b0 : n1519;
  /* TG68KdotC_Kernel.vhd:1257:25  */
  assign n1526 = clkena_lw ? n1525 : pcbase;
  /* TG68KdotC_Kernel.vhd:1255:25  */
  assign n1528 = reset ? 1'b1 : n1526;
  /* TG68KdotC_Kernel.vhd:1265:54  */
  assign n1529 = set[0]; // extract
  /* TG68KdotC_Kernel.vhd:1265:70  */
  assign n1530 = set[85]; // extract
  /* TG68KdotC_Kernel.vhd:1265:64  */
  assign n1531 = n1529 | n1530;
  /* TG68KdotC_Kernel.vhd:1266:58  */
  assign n1534 = set[3]; // extract
  /* TG68KdotC_Kernel.vhd:1266:73  */
  assign n1535 = set[86]; // extract
  /* TG68KdotC_Kernel.vhd:1266:67  */
  assign n1536 = n1534 | n1535;
  assign n1537 = set[88:87]; // extract
  /* TG68KdotC_Kernel.vhd:1268:52  */
  assign n1538 = set[47]; // extract
  /* TG68KdotC_Kernel.vhd:1268:67  */
  assign n1539 = set[48]; // extract
  /* TG68KdotC_Kernel.vhd:1268:61  */
  assign n1540 = n1538 | n1539;
  assign n1541 = set[84:49]; // extract
  assign n1542 = set[47:0]; // extract
  /* TG68KdotC_Kernel.vhd:1270:58  */
  assign n1543 = set_exec | set;
  /* TG68KdotC_Kernel.vhd:1271:67  */
  assign n1544 = set_exec[0]; // extract
  /* TG68KdotC_Kernel.vhd:1271:83  */
  assign n1545 = set[0]; // extract
  /* TG68KdotC_Kernel.vhd:1271:77  */
  assign n1546 = n1544 | n1545;
  /* TG68KdotC_Kernel.vhd:1271:99  */
  assign n1547 = set[85]; // extract
  /* TG68KdotC_Kernel.vhd:1271:93  */
  assign n1548 = n1546 | n1547;
  assign n1550 = n1543[84:0]; // extract
  /* TG68KdotC_Kernel.vhd:1272:71  */
  assign n1551 = set_exec[3]; // extract
  /* TG68KdotC_Kernel.vhd:1272:86  */
  assign n1552 = set[3]; // extract
  /* TG68KdotC_Kernel.vhd:1272:80  */
  assign n1553 = n1551 | n1552;
  /* TG68KdotC_Kernel.vhd:1272:101  */
  assign n1554 = set[86]; // extract
  /* TG68KdotC_Kernel.vhd:1272:95  */
  assign n1555 = n1553 | n1554;
  assign n1556 = n1543[88:87]; // extract
  /* TG68KdotC_Kernel.vhd:1269:33  */
  assign n1558 = setexecopc ? set_exec_tas : 1'b0;
  assign n1560 = {n1556, n1555, n1548, n1550};
  assign n1561 = {n1537, n1536, n1531, n1541, n1540, n1542};
  /* TG68KdotC_Kernel.vhd:1269:33  */
  assign n1562 = setexecopc ? n1560 : n1561;
  /* TG68KdotC_Kernel.vhd:1275:56  */
  assign n1563 = set[71]; // extract
  /* TG68KdotC_Kernel.vhd:1275:69  */
  assign n1564 = n1563 | setopcode;
  assign n1565 = n1562[88:72]; // extract
  assign n1566 = n1562[70:0]; // extract
  assign n1568 = {n1565, n1564, n1566};
  /* TG68KdotC_Kernel.vhd:1285:26  */
  assign n1576 = sndopc[11]; // extract
  /* TG68KdotC_Kernel.vhd:1286:48  */
  assign n1577 = reg_qa[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:1286:41  */
  assign n1579 = {1'b0, n1577};
  /* TG68KdotC_Kernel.vhd:1288:48  */
  assign n1580 = sndopc[10:6]; // extract
  /* TG68KdotC_Kernel.vhd:1288:41  */
  assign n1582 = {1'b0, n1580};
  /* TG68KdotC_Kernel.vhd:1285:17  */
  assign n1583 = n1576 ? n1579 : n1582;
  /* TG68KdotC_Kernel.vhd:1290:26  */
  assign n1584 = sndopc[11]; // extract
  /* TG68KdotC_Kernel.vhd:1294:61  */
  assign n1585 = sndopc[10:6]; // extract
  assign n1587 = n1586[31:5]; // extract
  assign n1588 = {n1587, n1585};
  /* TG68KdotC_Kernel.vhd:1290:17  */
  assign n1589 = n1584 ? reg_qa : n1588;
  /* TG68KdotC_Kernel.vhd:1298:26  */
  assign n1591 = sndopc[5]; // extract
  /* TG68KdotC_Kernel.vhd:1299:55  */
  assign n1592 = reg_qb[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:1299:67  */
  assign n1594 = n1592 - 5'b00001;
  /* TG68KdotC_Kernel.vhd:1301:55  */
  assign n1595 = sndopc[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:1301:67  */
  assign n1597 = n1595 - 5'b00001;
  /* TG68KdotC_Kernel.vhd:1298:17  */
  assign n1598 = n1591 ? n1594 : n1597;
  /* TG68KdotC_Kernel.vhd:1303:37  */
  assign n1599 = bf_width + bf_offset;
  /* TG68KdotC_Kernel.vhd:1304:43  */
  assign n1600 = bf_bhits[3]; // extract
  /* TG68KdotC_Kernel.vhd:1304:31  */
  assign n1601 = ~n1600;
  /* TG68KdotC_Kernel.vhd:1308:26  */
  assign n1602 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:1308:39  */
  assign n1604 = n1602 == 3'b111;
  /* TG68KdotC_Kernel.vhd:1309:41  */
  assign n1606 = 6'b100000 - bf_shift;
  /* TG68KdotC_Kernel.vhd:1308:17  */
  assign n1607 = n1604 ? n1606 : bf_shift;
  assign n1609 = n1607[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:1315:26  */
  assign n1610 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:1315:38  */
  assign n1612 = n1610 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1316:34  */
  assign n1613 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:1316:47  */
  assign n1615 = n1613 == 3'b111;
  /* TG68KdotC_Kernel.vhd:1317:53  */
  assign n1617 = bf_bhits + 6'b000001;
  /* TG68KdotC_Kernel.vhd:1319:47  */
  assign n1619 = 6'b011111 - bf_bhits;
  /* TG68KdotC_Kernel.vhd:1316:25  */
  assign n1620 = n1615 ? n1617 : n1619;
  assign n1622 = n1620[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:1323:34  */
  assign n1623 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:1323:47  */
  assign n1625 = n1623 == 3'b111;
  /* TG68KdotC_Kernel.vhd:1324:69  */
  assign n1626 = bf_bhits[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1324:60  */
  assign n1628 = {3'b000, n1626};
  /* TG68KdotC_Kernel.vhd:1324:53  */
  assign n1630 = 6'b011001 + n1628;
  assign n1632 = n1630[4:0]; // extract
  /* TG68KdotC_Kernel.vhd:1327:66  */
  assign n1633 = bf_bhits[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1327:57  */
  assign n1635 = 3'b111 - n1633;
  /* TG68KdotC_Kernel.vhd:1327:50  */
  assign n1637 = {3'b000, n1635};
  assign n1638 = {1'b0, n1632};
  /* TG68KdotC_Kernel.vhd:1323:25  */
  assign n1639 = n1625 ? n1638 : n1637;
  assign n1641 = n1583[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:1315:17  */
  assign n1642 = n1612 ? n1641 : 2'b00;
  assign n1643 = n1583[5]; // extract
  assign n1644 = n1583[2:0]; // extract
  assign n1645 = {1'b0, n1622};
  /* TG68KdotC_Kernel.vhd:1315:17  */
  assign n1646 = n1612 ? n1645 : n1639;
  /* TG68KdotC_Kernel.vhd:1332:30  */
  assign n1647 = bf_bhits[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1333:25  */
  assign n1649 = n1647 == 3'b000;
  /* TG68KdotC_Kernel.vhd:1335:25  */
  assign n1651 = n1647 == 3'b001;
  /* TG68KdotC_Kernel.vhd:1337:25  */
  assign n1653 = n1647 == 3'b010;
  /* TG68KdotC_Kernel.vhd:1339:25  */
  assign n1655 = n1647 == 3'b011;
  assign n1656 = {n1655, n1653, n1651, n1649};
  /* TG68KdotC_Kernel.vhd:1332:17  */
  always @*
    case (n1656)
      4'b1000: n1662 = 6'b100001;
      4'b0100: n1662 = 6'b100011;
      4'b0010: n1662 = 6'b100111;
      4'b0001: n1662 = 6'b101111;
      default: n1662 = 6'b100000;
    endcase
  /* TG68KdotC_Kernel.vhd:1344:28  */
  assign n1664 = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1344:17  */
  assign n1666 = n1664 ? 6'b100111 : n1662;
  /* TG68KdotC_Kernel.vhd:1354:24  */
  assign n1670 = exec[17]; // extract
  /* TG68KdotC_Kernel.vhd:1355:59  */
  assign n1671 = last_data_read[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:1355:41  */
  assign n1672 = flagssr & n1671;
  /* TG68KdotC_Kernel.vhd:1356:27  */
  assign n1673 = exec[18]; // extract
  /* TG68KdotC_Kernel.vhd:1357:59  */
  assign n1674 = last_data_read[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:1357:41  */
  assign n1675 = flagssr ^ n1674;
  /* TG68KdotC_Kernel.vhd:1358:27  */
  assign n1676 = exec[19]; // extract
  /* TG68KdotC_Kernel.vhd:1359:58  */
  assign n1677 = last_data_read[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:1359:41  */
  assign n1678 = flagssr | n1677;
  /* TG68KdotC_Kernel.vhd:1361:39  */
  assign n1679 = op2out[15:8]; // extract
  /* TG68KdotC_Kernel.vhd:1358:17  */
  assign n1680 = n1676 ? n1678 : n1679;
  /* TG68KdotC_Kernel.vhd:1356:17  */
  assign n1681 = n1673 ? n1675 : n1680;
  /* TG68KdotC_Kernel.vhd:1354:17  */
  assign n1682 = n1670 ? n1672 : n1681;
  /* TG68KdotC_Kernel.vhd:1373:62  */
  assign n1685 = flagssr[7]; // extract
  /* TG68KdotC_Kernel.vhd:1374:47  */
  assign n1686 = set[41]; // extract
  /* TG68KdotC_Kernel.vhd:1375:59  */
  assign n1687 = ~svmode;
  /* TG68KdotC_Kernel.vhd:1374:41  */
  assign n1688 = n1686 ? n1687 : presvmode;
  /* TG68KdotC_Kernel.vhd:1372:33  */
  assign n1689 = setopcode ? n1685 : make_trace;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1690 = n1759 ? n1688 : svmode;
  /* TG68KdotC_Kernel.vhd:1380:50  */
  assign n1691 = trap_berr | trap_illegal;
  /* TG68KdotC_Kernel.vhd:1380:70  */
  assign n1692 = n1691 | trap_addr_error;
  /* TG68KdotC_Kernel.vhd:1380:93  */
  assign n1693 = n1692 | trap_priv;
  /* TG68KdotC_Kernel.vhd:1380:110  */
  assign n1694 = n1693 | trap_1010;
  /* TG68KdotC_Kernel.vhd:1380:127  */
  assign n1695 = n1694 | trap_1111;
  assign n1697 = flagssr[7]; // extract
  /* TG68KdotC_Kernel.vhd:1380:33  */
  assign n1698 = n1695 ? 1'b0 : n1697;
  /* TG68KdotC_Kernel.vhd:1380:33  */
  assign n1700 = n1695 ? 1'b0 : n1689;
  /* TG68KdotC_Kernel.vhd:1384:39  */
  assign n1701 = set[41]; // extract
  /* TG68KdotC_Kernel.vhd:1385:54  */
  assign n1702 = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1386:55  */
  assign n1703 = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1387:50  */
  assign n1704 = ~presvmode;
  assign n1705 = n9425[2]; // extract
  /* TG68KdotC_Kernel.vhd:1384:33  */
  assign n1706 = n1701 ? n1704 : n1705;
  assign n1707 = flagssr[5]; // extract
  /* TG68KdotC_Kernel.vhd:1384:33  */
  assign n1708 = n1701 ? n1703 : n1707;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1709 = n1760 ? n1702 : presvmode;
  /* TG68KdotC_Kernel.vhd:1389:47  */
  assign n1711 = micro_state == 7'b0110110;
  /* TG68KdotC_Kernel.vhd:1389:33  */
  assign n1713 = n1711 ? 1'b0 : n1698;
  /* TG68KdotC_Kernel.vhd:1392:60  */
  assign n1715 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1392:51  */
  assign n1716 = n1715 & trap_trace;
  /* TG68KdotC_Kernel.vhd:1392:33  */
  assign n1718 = n1716 ? 1'b0 : n1700;
  /* TG68KdotC_Kernel.vhd:1395:40  */
  assign n1719 = exec[59]; // extract
  /* TG68KdotC_Kernel.vhd:1395:55  */
  assign n1720 = n1719 | set_stop;
  /* TG68KdotC_Kernel.vhd:1396:61  */
  assign n1721 = data_read[15:8]; // extract
  assign n1722 = flagssr[4:0]; // extract
  assign n1723 = flagssr[6]; // extract
  assign n1724 = {n1713, n1723, n1708, n1722};
  /* TG68KdotC_Kernel.vhd:1395:33  */
  assign n1725 = n1720 ? n1721 : n1724;
  /* TG68KdotC_Kernel.vhd:1398:50  */
  assign n1726 = trap_interrupt & interrupt;
  assign n1727 = n1725[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1398:33  */
  assign n1728 = n1726 ? ripl_nr : n1727;
  assign n1729 = n1725[7:3]; // extract
  /* TG68KdotC_Kernel.vhd:1401:40  */
  assign n1730 = exec[52]; // extract
  /* TG68KdotC_Kernel.vhd:1403:54  */
  assign n1731 = srin[5]; // extract
  /* TG68KdotC_Kernel.vhd:1404:43  */
  assign n1732 = exec[35]; // extract
  /* TG68KdotC_Kernel.vhd:1405:57  */
  assign n1733 = flagssr[5]; // extract
  /* TG68KdotC_Kernel.vhd:1404:33  */
  assign n1734 = n1732 ? n1733 : n1706;
  /* TG68KdotC_Kernel.vhd:1401:33  */
  assign n1735 = n1730 ? n1731 : n1734;
  assign n1736 = {n1729, n1728};
  /* TG68KdotC_Kernel.vhd:1401:33  */
  assign n1737 = n1730 ? srin : n1736;
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1739 = interrupt ? 1'b1 : n1735;
  /* TG68KdotC_Kernel.vhd:1410:39  */
  assign n1740 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:1410:42  */
  assign n1741 = ~n1740;
  assign n1744 = n1737[4]; // extract
  /* TG68KdotC_Kernel.vhd:1410:33  */
  assign n1745 = n1741 ? 1'b0 : n1744;
  assign n1746 = n1737[6]; // extract
  /* TG68KdotC_Kernel.vhd:1410:33  */
  assign n1747 = n1741 ? 1'b0 : n1746;
  assign n1750 = n1737[7]; // extract
  assign n1751 = n1737[5]; // extract
  assign n1753 = n1737[2:0]; // extract
  assign n1754 = n9425[2]; // extract
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1755 = clkena_lw ? n1739 : n1754;
  assign n1756 = {n1750, n1747, n1751, n1745, 1'b0, n1753};
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1757 = clkena_lw ? n1756 : flagssr;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1758 = clkena_lw ? n1718 : make_trace;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1759 = setopcode & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1760 = n1701 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1365:25  */
  assign n1761 = reset ? 1'b1 : n1755;
  /* TG68KdotC_Kernel.vhd:1365:25  */
  assign n1763 = reset ? 8'b00100111 : n1757;
  /* TG68KdotC_Kernel.vhd:1365:25  */
  assign n1765 = reset ? 1'b0 : n1758;
  /* TG68KdotC_Kernel.vhd:1365:25  */
  assign n1767 = reset ? 1'b1 : n1690;
  /* TG68KdotC_Kernel.vhd:1365:25  */
  assign n1769 = reset ? 1'b1 : n1709;
  /* TG68KdotC_Kernel.vhd:1447:39  */
  assign n1779 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:1489:27  */
  assign n1781 = rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1490:47  */
  assign n1783 = rot_cnt - 6'b000001;
  /* TG68KdotC_Kernel.vhd:1489:17  */
  assign n1785 = n1781 ? n1783 : 6'b000001;
  /* TG68KdotC_Kernel.vhd:1501:28  */
  assign n1791 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:1502:25  */
  assign n1793 = n1791 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1503:25  */
  assign n1795 = n1791 == 2'b01;
  assign n1796 = {n1795, n1793};
  /* TG68KdotC_Kernel.vhd:1501:17  */
  always @*
    case (n1796)
      2'b10: n1800 = 2'b01;
      2'b01: n1800 = 2'b00;
      default: n1800 = 2'b10;
    endcase
  /* TG68KdotC_Kernel.vhd:1507:32  */
  assign n1801 = exec_write_back & execopc;
  assign n1803 = n1788[83]; // extract
  /* TG68KdotC_Kernel.vhd:1507:17  */
  assign n1804 = n1801 ? 1'b1 : n1803;
  /* TG68KdotC_Kernel.vhd:1511:34  */
  assign n1807 = trap_berr & interrupt;
  /* TG68KdotC_Kernel.vhd:1513:37  */
  assign n1808 = ~presvmode;
  assign n1810 = n1788[41]; // extract
  /* TG68KdotC_Kernel.vhd:1511:17  */
  assign n1811 = n1817 ? 1'b1 : n1810;
  /* TG68KdotC_Kernel.vhd:1511:17  */
  assign n1814 = n1807 ? 2'b01 : 2'b00;
  /* TG68KdotC_Kernel.vhd:1511:17  */
  assign n1817 = n1808 & n1807;
  /* TG68KdotC_Kernel.vhd:1511:17  */
  assign n1822 = n1807 ? 7'b0110011 : 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1518:42  */
  assign n1824 = ~trapd;
  /* TG68KdotC_Kernel.vhd:1518:33  */
  assign n1825 = n1824 & trapmake;
  /* TG68KdotC_Kernel.vhd:1519:31  */
  assign n1826 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:1519:59  */
  assign n1827 = trap_trapv | set_z_error;
  /* TG68KdotC_Kernel.vhd:1519:85  */
  assign n1828 = exec[43]; // extract
  /* TG68KdotC_Kernel.vhd:1519:78  */
  assign n1829 = n1827 | n1828;
  /* TG68KdotC_Kernel.vhd:1519:39  */
  assign n1830 = n1829 & n1826;
  /* TG68KdotC_Kernel.vhd:1519:25  */
  assign n1833 = n1830 ? 7'b0110010 : 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1524:46  */
  assign n1834 = ~use_vbr_stackframe;
  assign n1836 = n1788[25]; // extract
  /* TG68KdotC_Kernel.vhd:1518:17  */
  assign n1837 = n1844 ? 1'b1 : n1836;
  /* TG68KdotC_Kernel.vhd:1528:37  */
  assign n1838 = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1518:17  */
  assign n1840 = n1845 ? 1'b1 : n1811;
  /* TG68KdotC_Kernel.vhd:1518:17  */
  assign n1842 = n1825 ? 2'b01 : n1814;
  /* TG68KdotC_Kernel.vhd:1518:17  */
  assign n1844 = n1834 & n1825;
  /* TG68KdotC_Kernel.vhd:1518:17  */
  assign n1845 = n1838 & n1825;
  /* TG68KdotC_Kernel.vhd:1518:17  */
  assign n1848 = n1825 ? n1833 : n1822;
  /* TG68KdotC_Kernel.vhd:1533:31  */
  assign n1850 = micro_state == 7'b0100111;
  /* TG68KdotC_Kernel.vhd:1533:55  */
  assign n1851 = trap_trace & interrupt;
  /* TG68KdotC_Kernel.vhd:1533:37  */
  assign n1852 = n1850 | n1851;
  /* TG68KdotC_Kernel.vhd:1535:50  */
  assign n1853 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:1535:43  */
  assign n1854 = n1853 & trap_trace;
  /* TG68KdotC_Kernel.vhd:1535:25  */
  assign n1857 = n1854 ? 7'b0110010 : 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1545:37  */
  assign n1858 = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1533:17  */
  assign n1860 = n1863 ? 1'b1 : n1840;
  /* TG68KdotC_Kernel.vhd:1533:17  */
  assign n1862 = n1852 ? 2'b01 : n1842;
  /* TG68KdotC_Kernel.vhd:1533:17  */
  assign n1863 = n1858 & n1852;
  /* TG68KdotC_Kernel.vhd:1533:17  */
  assign n1864 = n1852 ? n1857 : n1848;
  /* TG68KdotC_Kernel.vhd:1550:24  */
  assign n1866 = micro_state == 7'b0100111;
  /* TG68KdotC_Kernel.vhd:1550:51  */
  assign n1867 = trap_trace & interrupt;
  /* TG68KdotC_Kernel.vhd:1550:31  */
  assign n1868 = n1866 | n1867;
  /* TG68KdotC_Kernel.vhd:1551:24  */
  assign n1869 = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1550:9  */
  assign n1871 = n1874 ? 1'b1 : n1860;
  /* TG68KdotC_Kernel.vhd:1550:9  */
  assign n1873 = n1868 ? 2'b01 : n1862;
  /* TG68KdotC_Kernel.vhd:1550:9  */
  assign n1874 = n1869 & n1868;
  /* TG68KdotC_Kernel.vhd:1557:46  */
  assign n1875 = flagssr[5]; // extract
  /* TG68KdotC_Kernel.vhd:1557:49  */
  assign n1876 = n1875 != presvmode;
  /* TG68KdotC_Kernel.vhd:1557:35  */
  assign n1877 = n1876 & setexecopc;
  /* TG68KdotC_Kernel.vhd:1557:17  */
  assign n1879 = n1877 ? 1'b1 : n1871;
  /* TG68KdotC_Kernel.vhd:1563:34  */
  assign n1880 = trap_interrupt & interrupt;
  /* TG68KdotC_Kernel.vhd:1563:17  */
  assign n1883 = n1880 ? 2'b10 : n1873;
  /* TG68KdotC_Kernel.vhd:1563:17  */
  assign n1884 = n1880 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1563:17  */
  assign n1886 = n1880 ? 7'b0100111 : n1864;
  /* TG68KdotC_Kernel.vhd:1570:23  */
  assign n1887 = set[41]; // extract
  /* TG68KdotC_Kernel.vhd:1570:17  */
  assign n1892 = n1887 ? 1'b1 : 1'b0;
  assign n1894 = {1'b1, 1'b1};
  assign n1895 = n1788[66:65]; // extract
  /* TG68KdotC_Kernel.vhd:1570:17  */
  assign n1896 = n1887 ? n1894 : n1895;
  /* TG68KdotC_Kernel.vhd:1576:27  */
  assign n1899 = ~ea_only;
  /* TG68KdotC_Kernel.vhd:1576:39  */
  assign n1900 = set[62]; // extract
  /* TG68KdotC_Kernel.vhd:1576:32  */
  assign n1901 = n1900 & n1899;
  /* TG68KdotC_Kernel.vhd:1576:17  */
  assign n1903 = n1901 ? 2'b10 : n1883;
  /* TG68KdotC_Kernel.vhd:1582:28  */
  assign n1904 = setstate[1]; // extract
  /* TG68KdotC_Kernel.vhd:1582:52  */
  assign n1905 = set_datatype[1]; // extract
  /* TG68KdotC_Kernel.vhd:1582:36  */
  assign n1906 = n1905 & n1904;
  assign n1908 = n1788[73]; // extract
  /* TG68KdotC_Kernel.vhd:1582:17  */
  assign n1909 = n1906 ? 1'b1 : n1908;
  /* TG68KdotC_Kernel.vhd:1586:38  */
  assign n1912 = decodeopc & ea_build_now;
  /* TG68KdotC_Kernel.vhd:1586:64  */
  assign n1913 = exec[42]; // extract
  /* TG68KdotC_Kernel.vhd:1586:57  */
  assign n1914 = n1912 | n1913;
  /* TG68KdotC_Kernel.vhd:1587:36  */
  assign n1915 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1591:50  */
  assign n1917 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:1593:58  */
  assign n1919 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1593:70  */
  assign n1921 = n1919 == 3'b111;
  assign n1923 = n1788[50]; // extract
  /* TG68KdotC_Kernel.vhd:1591:41  */
  assign n1924 = n1928 ? 1'b1 : n1923;
  assign n1925 = n1788[46]; // extract
  /* TG68KdotC_Kernel.vhd:1591:41  */
  assign n1926 = n1917 ? 1'b1 : n1925;
  /* TG68KdotC_Kernel.vhd:1591:41  */
  assign n1928 = n1921 & n1917;
  /* TG68KdotC_Kernel.vhd:1597:50  */
  assign n1929 = opcode[5]; // extract
  /* TG68KdotC_Kernel.vhd:1599:58  */
  assign n1931 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1599:70  */
  assign n1933 = n1931 == 3'b111;
  /* TG68KdotC_Kernel.vhd:1597:41  */
  assign n1935 = n1938 ? 1'b1 : n1924;
  assign n1936 = n1788[47]; // extract
  /* TG68KdotC_Kernel.vhd:1597:41  */
  assign n1937 = n1929 ? 1'b1 : n1936;
  /* TG68KdotC_Kernel.vhd:1597:41  */
  assign n1938 = n1933 & n1929;
  /* TG68KdotC_Kernel.vhd:1588:33  */
  assign n1940 = n1915 == 3'b010;
  /* TG68KdotC_Kernel.vhd:1588:43  */
  assign n1942 = n1915 == 3'b011;
  /* TG68KdotC_Kernel.vhd:1588:43  */
  assign n1943 = n1940 | n1942;
  /* TG68KdotC_Kernel.vhd:1588:49  */
  assign n1945 = n1915 == 3'b100;
  /* TG68KdotC_Kernel.vhd:1588:49  */
  assign n1946 = n1943 | n1945;
  /* TG68KdotC_Kernel.vhd:1603:33  */
  assign n1948 = n1915 == 3'b101;
  /* TG68KdotC_Kernel.vhd:1605:33  */
  assign n1950 = n1915 == 3'b110;
  /* TG68KdotC_Kernel.vhd:1609:52  */
  assign n1951 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1610:49  */
  assign n1953 = n1951 == 3'b000;
  /* TG68KdotC_Kernel.vhd:1612:49  */
  assign n1956 = n1951 == 3'b001;
  /* TG68KdotC_Kernel.vhd:1615:49  */
  assign n1959 = n1951 == 3'b010;
  /* TG68KdotC_Kernel.vhd:1620:49  */
  assign n1962 = n1951 == 3'b011;
  /* TG68KdotC_Kernel.vhd:1629:68  */
  assign n1964 = datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:1629:57  */
  assign n1966 = n1964 ? 1'b1 : n1909;
  /* TG68KdotC_Kernel.vhd:1626:49  */
  assign n1968 = n1951 == 3'b100;
  assign n1969 = {n1968, n1962, n1959, n1956, n1953};
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1972 = 1'b1;
      5'b01000: n1972 = 1'b0;
      5'b00100: n1972 = 1'b0;
      5'b00010: n1972 = 1'b0;
      5'b00001: n1972 = 1'b0;
      default: n1972 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1975 = 1'b0;
      5'b01000: n1975 = 1'b1;
      5'b00100: n1975 = 1'b0;
      5'b00010: n1975 = 1'b0;
      5'b00001: n1975 = 1'b0;
      default: n1975 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1978 = 1'b1;
      5'b01000: n1978 = 1'b0;
      5'b00100: n1978 = 1'b0;
      5'b00010: n1978 = 1'b0;
      5'b00001: n1978 = 1'b0;
      default: n1978 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1982 = 1'b0;
      5'b01000: n1982 = 1'b1;
      5'b00100: n1982 = 1'b1;
      5'b00010: n1982 = 1'b0;
      5'b00001: n1982 = 1'b0;
      default: n1982 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1986 = 1'b0;
      5'b01000: n1986 = 1'b1;
      5'b00100: n1986 = 1'b1;
      5'b00010: n1986 = 1'b0;
      5'b00001: n1986 = 1'b0;
      default: n1986 = 1'b0;
    endcase
  assign n1987 = n1788[22]; // extract
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1988 = n1987;
      5'b01000: n1988 = 1'b1;
      5'b00100: n1988 = 1'b1;
      5'b00010: n1988 = n1987;
      5'b00001: n1988 = n1987;
      default: n1988 = n1987;
    endcase
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1989 = n1966;
      5'b01000: n1989 = n1909;
      5'b00100: n1989 = n1909;
      5'b00010: n1989 = 1'b1;
      5'b00001: n1989 = n1909;
      default: n1989 = n1909;
    endcase
  /* TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n1969)
      5'b10000: n1994 = n1886;
      5'b01000: n1994 = 7'b0000101;
      5'b00100: n1994 = 7'b0000100;
      5'b00010: n1994 = 7'b0000010;
      5'b00001: n1994 = 7'b0000010;
      default: n1994 = n1886;
    endcase
  /* TG68KdotC_Kernel.vhd:1608:33  */
  assign n1996 = n1915 == 3'b111;
  assign n1997 = {n1996, n1950, n1948, n1946};
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2000 = n1972;
      4'b0100: n2000 = 1'b0;
      4'b0010: n2000 = 1'b0;
      4'b0001: n2000 = 1'b1;
      default: n2000 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2003 = n1975;
      4'b0100: n2003 = 1'b1;
      4'b0010: n2003 = 1'b0;
      4'b0001: n2003 = 1'b0;
      default: n2003 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2005 = n1978;
      4'b0100: n2005 = 1'b0;
      4'b0010: n2005 = 1'b0;
      4'b0001: n2005 = 1'b0;
      default: n2005 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2007 = n1982;
      4'b0100: n2007 = 1'b0;
      4'b0010: n2007 = 1'b0;
      4'b0001: n2007 = 1'b0;
      default: n2007 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2009 = n1986;
      4'b0100: n2009 = 1'b0;
      4'b0010: n2009 = 1'b0;
      4'b0001: n2009 = 1'b0;
      default: n2009 = 1'b0;
    endcase
  assign n2010 = n1788[22]; // extract
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2011 = n1988;
      4'b0100: n2011 = n2010;
      4'b0010: n2011 = n2010;
      4'b0001: n2011 = n2010;
      default: n2011 = n2010;
    endcase
  assign n2012 = n1788[46]; // extract
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2013 = n2012;
      4'b0100: n2013 = n2012;
      4'b0010: n2013 = n2012;
      4'b0001: n2013 = n1926;
      default: n2013 = n2012;
    endcase
  assign n2014 = n1788[47]; // extract
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2015 = n2014;
      4'b0100: n2015 = n2014;
      4'b0010: n2015 = n2014;
      4'b0001: n2015 = n1937;
      default: n2015 = n2014;
    endcase
  assign n2016 = n1788[50]; // extract
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2017 = n2016;
      4'b0100: n2017 = n2016;
      4'b0010: n2017 = n2016;
      4'b0001: n2017 = n1935;
      default: n2017 = n2016;
    endcase
  assign n2018 = n1788[62]; // extract
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2019 = n2018;
      4'b0100: n2019 = n2018;
      4'b0010: n2019 = n2018;
      4'b0001: n2019 = 1'b1;
      default: n2019 = n2018;
    endcase
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2020 = n1989;
      4'b0100: n2020 = n1909;
      4'b0010: n2020 = n1909;
      4'b0001: n2020 = n1909;
      default: n2020 = n1909;
    endcase
  /* TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n1997)
      4'b1000: n2023 = n1994;
      4'b0100: n2023 = 7'b0000101;
      4'b0010: n2023 = 7'b0000100;
      4'b0001: n2023 = n1886;
      default: n2023 = n1886;
    endcase
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2025 = n1914 ? n2000 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2028 = n1914 ? n2003 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2031 = n1914 ? n2005 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2034 = n1914 ? n2007 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2037 = n1914 ? n2009 : 1'b0;
  assign n2039 = {n2015, n2013};
  assign n2040 = n1788[22]; // extract
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2041 = n1914 ? n2011 : n2040;
  assign n2042 = n1788[47:46]; // extract
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2043 = n1914 ? n2039 : n2042;
  assign n2044 = n1788[50]; // extract
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2045 = n1914 ? n2017 : n2044;
  assign n2046 = n1788[62]; // extract
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2047 = n1914 ? n2019 : n2046;
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2048 = n1914 ? n2020 : n1909;
  assign n2054 = n1788[49:48]; // extract
  assign n2055 = n1788[64:63]; // extract
  /* TG68KdotC_Kernel.vhd:1586:17  */
  assign n2057 = n1914 ? n2023 : n1886;
  /* TG68KdotC_Kernel.vhd:1640:28  */
  assign n2058 = opcode[15:12]; // extract
  /* TG68KdotC_Kernel.vhd:1643:34  */
  assign n2059 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:1643:52  */
  assign n2060 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1643:64  */
  assign n2062 = n2060 == 3'b001;
  /* TG68KdotC_Kernel.vhd:1643:42  */
  assign n2063 = n2062 & n2059;
  /* TG68KdotC_Kernel.vhd:1647:42  */
  assign n2066 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1647:45  */
  assign n2067 = ~n2066;
  assign n2071 = n1788[37]; // extract
  /* TG68KdotC_Kernel.vhd:1647:33  */
  assign n2072 = n2067 ? 1'b1 : n2071;
  /* TG68KdotC_Kernel.vhd:1647:33  */
  assign n2074 = n2067 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1647:33  */
  assign n2076 = n2067 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1653:50  */
  assign n2077 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:1652:33  */
  assign n2079 = n2085 ? 1'b1 : n2072;
  /* TG68KdotC_Kernel.vhd:1656:50  */
  assign n2080 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1656:53  */
  assign n2081 = ~n2080;
  /* TG68KdotC_Kernel.vhd:1652:33  */
  assign n2083 = n2084 ? 1'b1 : n2031;
  /* TG68KdotC_Kernel.vhd:1652:33  */
  assign n2084 = n2081 & decodeopc;
  /* TG68KdotC_Kernel.vhd:1652:33  */
  assign n2085 = n2077 & decodeopc;
  /* TG68KdotC_Kernel.vhd:1652:33  */
  assign n2087 = decodeopc ? 7'b1001010 : n2057;
  /* TG68KdotC_Kernel.vhd:1661:33  */
  assign n2090 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1665:42  */
  assign n2091 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:1665:59  */
  assign n2092 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1665:72  */
  assign n2094 = n2092 == 3'b100;
  /* TG68KdotC_Kernel.vhd:1665:50  */
  assign n2095 = n2091 | n2094;
  /* TG68KdotC_Kernel.vhd:1666:50  */
  assign n2096 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1666:62  */
  assign n2098 = n2096 != 3'b001;
  /* TG68KdotC_Kernel.vhd:1667:51  */
  assign n2099 = opcode[8:3]; // extract
  /* TG68KdotC_Kernel.vhd:1667:63  */
  assign n2101 = n2099 != 6'b000111;
  /* TG68KdotC_Kernel.vhd:1667:83  */
  assign n2102 = opcode[2]; // extract
  /* TG68KdotC_Kernel.vhd:1667:86  */
  assign n2103 = ~n2102;
  /* TG68KdotC_Kernel.vhd:1667:74  */
  assign n2104 = n2101 | n2103;
  /* TG68KdotC_Kernel.vhd:1666:70  */
  assign n2105 = n2104 & n2098;
  /* TG68KdotC_Kernel.vhd:1668:51  */
  assign n2106 = opcode[8:2]; // extract
  /* TG68KdotC_Kernel.vhd:1668:63  */
  assign n2108 = n2106 != 7'b1001111;
  /* TG68KdotC_Kernel.vhd:1668:84  */
  assign n2109 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:1668:96  */
  assign n2111 = n2109 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1668:75  */
  assign n2112 = n2108 | n2111;
  /* TG68KdotC_Kernel.vhd:1667:92  */
  assign n2113 = n2112 & n2105;
  /* TG68KdotC_Kernel.vhd:1669:51  */
  assign n2114 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:1669:63  */
  assign n2116 = n2114 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1669:78  */
  assign n2117 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1669:90  */
  assign n2119 = n2117 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1669:69  */
  assign n2120 = n2116 | n2119;
  /* TG68KdotC_Kernel.vhd:1669:107  */
  assign n2121 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1669:119  */
  assign n2123 = n2121 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1669:98  */
  assign n2124 = n2120 | n2123;
  /* TG68KdotC_Kernel.vhd:1668:103  */
  assign n2125 = n2124 & n2113;
  /* TG68KdotC_Kernel.vhd:1672:58  */
  assign n2128 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:1672:70  */
  assign n2130 = n2128 != 2'b00;
  /* TG68KdotC_Kernel.vhd:1673:66  */
  assign n2131 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1673:78  */
  assign n2133 = n2131 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1673:57  */
  assign n2136 = n2133 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1672:49  */
  assign n2139 = n2130 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1672:49  */
  assign n2141 = n2130 ? n2136 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1678:58  */
  assign n2142 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1678:70  */
  assign n2144 = n2142 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1678:49  */
  assign n2147 = n2144 ? 2'b10 : 2'b00;
  /* TG68KdotC_Kernel.vhd:1683:58  */
  assign n2148 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:1683:61  */
  assign n2149 = ~n2148;
  assign n2152 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2153 = n2178 ? 1'b1 : n2152;
  assign n2154 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2155 = n2180 ? 1'b1 : n2154;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2157 = n2187 ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:1683:49  */
  assign n2160 = n2149 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1683:49  */
  assign n2162 = decodeopc & n2149;
  /* TG68KdotC_Kernel.vhd:1683:49  */
  assign n2164 = decodeopc & n2149;
  /* TG68KdotC_Kernel.vhd:1683:49  */
  assign n2165 = decodeopc & n2149;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2166 = n2125 ? n2147 : n1800;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2168 = n2125 ? n2139 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2171 = n2125 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2174 = n2125 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2176 = n2125 ? n2160 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2178 = n2162 & n2125;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2180 = n2164 & n2125;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2182 = n2125 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2184 = n2125 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2186 = n2125 ? n2141 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1666:41  */
  assign n2187 = n2165 & n2125;
  /* TG68KdotC_Kernel.vhd:1696:45  */
  assign n2188 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:1696:57  */
  assign n2190 = n2188 == 3'b011;
  /* TG68KdotC_Kernel.vhd:1697:47  */
  assign n2191 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:1698:58  */
  assign n2192 = opcode[11]; // extract
  /* TG68KdotC_Kernel.vhd:1699:67  */
  assign n2193 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:1699:80  */
  assign n2195 = n2193 != 2'b00;
  /* TG68KdotC_Kernel.vhd:1700:66  */
  assign n2196 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1700:78  */
  assign n2198 = n2196 != 2'b00;
  /* TG68KdotC_Kernel.vhd:1699:87  */
  assign n2199 = n2198 & n2195;
  /* TG68KdotC_Kernel.vhd:1700:96  */
  assign n2200 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1700:108  */
  assign n2202 = n2200 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1700:125  */
  assign n2203 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1700:137  */
  assign n2205 = n2203 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1700:116  */
  assign n2206 = n2202 | n2205;
  /* TG68KdotC_Kernel.vhd:1700:85  */
  assign n2207 = n2206 & n2199;
  /* TG68KdotC_Kernel.vhd:1701:67  */
  assign n2208 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:1701:86  */
  assign n2209 = opcode[5:0]; // extract
  /* TG68KdotC_Kernel.vhd:1701:98  */
  assign n2211 = n2209 == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1701:76  */
  assign n2212 = n2211 & n2208;
  /* TG68KdotC_Kernel.vhd:1700:145  */
  assign n2213 = n2207 | n2212;
  /* TG68KdotC_Kernel.vhd:1702:76  */
  assign n2214 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:1703:73  */
  assign n2216 = n2214 == 2'b01;
  /* TG68KdotC_Kernel.vhd:1704:73  */
  assign n2218 = n2214 == 2'b10;
  assign n2219 = {n2218, n2216};
  /* TG68KdotC_Kernel.vhd:1702:65  */
  always @*
    case (n2219)
      2'b10: n2223 = 2'b01;
      2'b01: n2223 = 2'b00;
      default: n2223 = 2'b10;
    endcase
  /* TG68KdotC_Kernel.vhd:1707:74  */
  assign n2224 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:1707:93  */
  assign n2225 = opcode[5:0]; // extract
  /* TG68KdotC_Kernel.vhd:1707:105  */
  assign n2227 = n2225 == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1707:83  */
  assign n2228 = n2227 & n2224;
  assign n2230 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1708:73  */
  assign n2231 = decodeopc ? 1'b1 : n2230;
  /* TG68KdotC_Kernel.vhd:1708:73  */
  assign n2233 = decodeopc ? 7'b0111001 : n2057;
  assign n2236 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1713:73  */
  assign n2237 = decodeopc ? 1'b1 : n2236;
  assign n2238 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1713:73  */
  assign n2239 = decodeopc ? 1'b1 : n2238;
  /* TG68KdotC_Kernel.vhd:1713:73  */
  assign n2241 = decodeopc ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:1718:87  */
  assign n2243 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1718:93  */
  assign n2244 = nextpass & n2243;
  /* TG68KdotC_Kernel.vhd:1718:73  */
  assign n2250 = n2244 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:1718:73  */
  assign n2253 = n2244 ? 1'b1 : 1'b0;
  assign n2254 = n1788[26]; // extract
  /* TG68KdotC_Kernel.vhd:1718:73  */
  assign n2255 = n2244 ? 1'b1 : n2254;
  assign n2256 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1718:73  */
  assign n2257 = n2244 ? 1'b1 : n2256;
  assign n2258 = n1788[84]; // extract
  /* TG68KdotC_Kernel.vhd:1718:73  */
  assign n2259 = n2244 ? 1'b1 : n2258;
  assign n2260 = n1788[86]; // extract
  /* TG68KdotC_Kernel.vhd:1718:73  */
  assign n2261 = n2244 ? 1'b1 : n2260;
  /* TG68KdotC_Kernel.vhd:1718:73  */
  assign n2263 = n2244 ? 7'b0110111 : n2241;
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2264 = n2228 ? n1903 : n2250;
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2266 = n2228 ? 1'b0 : n2253;
  assign n2267 = n1788[26]; // extract
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2268 = n2228 ? n2267 : n2255;
  assign n2269 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2270 = n2228 ? n2269 : n2237;
  assign n2271 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2272 = n2228 ? n2271 : n2257;
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2273 = n2228 ? n2231 : n2239;
  assign n2274 = n1788[84]; // extract
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2275 = n2228 ? n2274 : n2259;
  assign n2276 = n1788[86]; // extract
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2277 = n2228 ? n2276 : n2261;
  /* TG68KdotC_Kernel.vhd:1707:65  */
  assign n2278 = n2228 ? n2233 : n2263;
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2279 = n2213 ? n2223 : n1800;
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2280 = n2213 ? n2264 : n1903;
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2282 = n2213 ? n2266 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2285 = n2213 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2288 = n2213 ? 1'b0 : 1'b1;
  assign n2289 = n1788[26]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2290 = n2868 ? n2268 : n2289;
  assign n2291 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2292 = n2213 ? n2270 : n2291;
  assign n2293 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2294 = n2397 ? n2272 : n2293;
  assign n2295 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2296 = n2213 ? n2273 : n2295;
  assign n2297 = n1788[84]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2298 = n2890 ? n2275 : n2297;
  assign n2299 = n1788[86]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2300 = n2892 ? n2277 : n2299;
  /* TG68KdotC_Kernel.vhd:1699:57  */
  assign n2301 = n2213 ? n2278 : n2057;
  /* TG68KdotC_Kernel.vhd:1733:66  */
  assign n2302 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:1733:79  */
  assign n2304 = n2302 != 2'b11;
  /* TG68KdotC_Kernel.vhd:1734:66  */
  assign n2305 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1734:78  */
  assign n2307 = n2305 != 2'b00;
  /* TG68KdotC_Kernel.vhd:1733:86  */
  assign n2308 = n2307 & n2304;
  /* TG68KdotC_Kernel.vhd:1734:95  */
  assign n2309 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1734:107  */
  assign n2311 = n2309 != 3'b011;
  /* TG68KdotC_Kernel.vhd:1734:85  */
  assign n2312 = n2311 & n2308;
  /* TG68KdotC_Kernel.vhd:1734:125  */
  assign n2313 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1734:137  */
  assign n2315 = n2313 != 3'b100;
  /* TG68KdotC_Kernel.vhd:1734:115  */
  assign n2316 = n2315 & n2312;
  /* TG68KdotC_Kernel.vhd:1734:155  */
  assign n2317 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:1734:167  */
  assign n2319 = n2317 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1734:145  */
  assign n2320 = n2319 & n2316;
  /* TG68KdotC_Kernel.vhd:1736:83  */
  assign n2322 = opcode[10:9]; // extract
  assign n2325 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1737:65  */
  assign n2326 = decodeopc ? 1'b1 : n2325;
  assign n2327 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2328 = n2373 ? 1'b1 : n2327;
  /* TG68KdotC_Kernel.vhd:1737:65  */
  assign n2330 = decodeopc ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:1742:71  */
  assign n2331 = set[62]; // extract
  assign n2334 = n1788[39]; // extract
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2335 = n2367 ? 1'b1 : n2334;
  assign n2336 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2337 = n2371 ? 1'b1 : n2336;
  /* TG68KdotC_Kernel.vhd:1746:79  */
  assign n2339 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1746:85  */
  assign n2340 = nextpass & n2339;
  /* TG68KdotC_Kernel.vhd:1749:88  */
  assign n2343 = exe_datatype != 2'b00;
  /* TG68KdotC_Kernel.vhd:1749:73  */
  assign n2346 = n2343 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2348 = n2356 ? 2'b10 : n1903;
  /* TG68KdotC_Kernel.vhd:1746:65  */
  assign n2350 = n2340 ? n2346 : 1'b0;
  assign n2351 = n1788[82]; // extract
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2352 = n2375 ? 1'b1 : n2351;
  /* TG68KdotC_Kernel.vhd:1746:65  */
  assign n2354 = n2340 ? 7'b1000001 : n2330;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2355 = n2320 ? n2322 : n1800;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2356 = n2340 & n2320;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2359 = n2320 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2362 = n2320 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2364 = n2320 ? n2350 : 1'b0;
  assign n2365 = {1'b1, n2326};
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2367 = n2331 & n2320;
  assign n2368 = n1788[43:42]; // extract
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2369 = n2320 ? n2365 : n2368;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2371 = n2331 & n2320;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2373 = decodeopc & n2320;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2375 = n2340 & n2320;
  /* TG68KdotC_Kernel.vhd:1733:57  */
  assign n2376 = n2320 ? n2354 : n2057;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2377 = n2192 ? n2279 : n2355;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2378 = n2192 ? n2280 : n2348;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2380 = n2192 ? n2282 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2381 = n2192 ? n2285 : n2359;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2382 = n2192 ? n2288 : n2362;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2384 = n2192 ? 1'b0 : n2364;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2386 = n2213 & n2192;
  assign n2387 = n1788[39]; // extract
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2388 = n2192 ? n2387 : n2335;
  assign n2389 = n2369[0]; // extract
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2390 = n2192 ? n2292 : n2389;
  assign n2391 = n2369[1]; // extract
  assign n2392 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2393 = n2192 ? n2392 : n2391;
  assign n2394 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2395 = n2192 ? n2394 : n2337;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2397 = n2213 & n2192;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2398 = n2192 ? n2296 : n2328;
  assign n2399 = n1788[82]; // extract
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2400 = n2192 ? n2399 : n2352;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2402 = n2213 & n2192;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2404 = n2213 & n2192;
  /* TG68KdotC_Kernel.vhd:1698:49  */
  assign n2405 = n2192 ? n2301 : n2376;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2406 = n2852 ? n2377 : n1800;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2407 = n2191 ? n2378 : n1903;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2409 = n2191 ? n2380 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2411 = n2191 ? n2381 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2413 = n2191 ? n2382 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2415 = n2191 ? n2384 : 1'b0;
  assign n2416 = {n2393, n2390};
  assign n2417 = {n2294, n2395};
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2419 = n2386 & n2191;
  assign n2420 = n1788[39]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2421 = n2870 ? n2388 : n2420;
  assign n2422 = n1788[43:42]; // extract
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2423 = n2191 ? n2416 : n2422;
  assign n2424 = n1788[56:55]; // extract
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2425 = n2191 ? n2417 : n2424;
  assign n2426 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2427 = n2191 ? n2398 : n2426;
  assign n2428 = n1788[82]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2429 = n2888 ? n2400 : n2428;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2431 = n2402 & n2191;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2433 = n2404 & n2191;
  /* TG68KdotC_Kernel.vhd:1697:41  */
  assign n2434 = n2191 ? n2405 : n2057;
  /* TG68KdotC_Kernel.vhd:1763:45  */
  assign n2435 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1763:58  */
  assign n2437 = n2435 == 3'b111;
  /* TG68KdotC_Kernel.vhd:1764:47  */
  assign n2438 = CPU[0]; // extract
  /* TG68KdotC_Kernel.vhd:1764:65  */
  assign n2439 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:1764:77  */
  assign n2441 = n2439 != 2'b11;
  /* TG68KdotC_Kernel.vhd:1764:55  */
  assign n2442 = n2441 & n2438;
  /* TG68KdotC_Kernel.vhd:1764:94  */
  assign n2443 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1764:106  */
  assign n2445 = n2443 != 2'b00;
  /* TG68KdotC_Kernel.vhd:1764:84  */
  assign n2446 = n2445 & n2442;
  /* TG68KdotC_Kernel.vhd:1764:124  */
  assign n2447 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1764:136  */
  assign n2449 = n2447 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1764:153  */
  assign n2450 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1764:165  */
  assign n2452 = n2450 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1764:144  */
  assign n2453 = n2449 | n2452;
  /* TG68KdotC_Kernel.vhd:1764:113  */
  assign n2454 = n2453 & n2446;
  /* TG68KdotC_Kernel.vhd:1765:49  */
  assign n2457 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1765:49  */
  assign n2460 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1764:41  */
  assign n2462 = n2454 ? n2457 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1764:41  */
  assign n2464 = n2454 ? n2460 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:50  */
  assign n2465 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:1778:62  */
  assign n2467 = n2465 != 2'b11;
  /* TG68KdotC_Kernel.vhd:1778:79  */
  assign n2468 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1778:91  */
  assign n2470 = n2468 != 3'b001;
  /* TG68KdotC_Kernel.vhd:1778:69  */
  assign n2471 = n2470 & n2467;
  /* TG68KdotC_Kernel.vhd:1779:58  */
  assign n2472 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1779:71  */
  assign n2474 = n2472 == 3'b000;
  /* TG68KdotC_Kernel.vhd:1780:66  */
  assign n2475 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1780:78  */
  assign n2477 = n2475 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1780:95  */
  assign n2478 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1780:107  */
  assign n2480 = n2478 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1780:86  */
  assign n2481 = n2477 | n2480;
  /* TG68KdotC_Kernel.vhd:1780:123  */
  assign n2482 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1780:135  */
  assign n2484 = n2482 == 3'b100;
  /* TG68KdotC_Kernel.vhd:1780:152  */
  assign n2485 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1780:155  */
  assign n2486 = ~n2485;
  /* TG68KdotC_Kernel.vhd:1780:142  */
  assign n2487 = n2486 & n2484;
  /* TG68KdotC_Kernel.vhd:1780:113  */
  assign n2488 = n2481 | n2487;
  /* TG68KdotC_Kernel.vhd:1780:57  */
  assign n2492 = n2488 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1780:57  */
  assign n2495 = n2488 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1780:57  */
  assign n2497 = n2488 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1779:49  */
  assign n2499 = n2474 ? n2492 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1779:49  */
  assign n2501 = n2474 ? n2495 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1779:49  */
  assign n2503 = n2474 ? n2497 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1787:58  */
  assign n2504 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1787:71  */
  assign n2506 = n2504 == 3'b001;
  /* TG68KdotC_Kernel.vhd:1788:66  */
  assign n2507 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1788:78  */
  assign n2509 = n2507 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1788:95  */
  assign n2510 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1788:107  */
  assign n2512 = n2510 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1788:86  */
  assign n2513 = n2509 | n2512;
  /* TG68KdotC_Kernel.vhd:1788:123  */
  assign n2514 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1788:135  */
  assign n2516 = n2514 == 3'b100;
  /* TG68KdotC_Kernel.vhd:1788:152  */
  assign n2517 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1788:155  */
  assign n2518 = ~n2517;
  /* TG68KdotC_Kernel.vhd:1788:142  */
  assign n2519 = n2518 & n2516;
  /* TG68KdotC_Kernel.vhd:1788:113  */
  assign n2520 = n2513 | n2519;
  /* TG68KdotC_Kernel.vhd:1788:57  */
  assign n2523 = n2520 ? n2499 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1788:57  */
  assign n2525 = n2520 ? n2501 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1788:57  */
  assign n2527 = n2520 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1787:49  */
  assign n2528 = n2506 ? n2523 : n2499;
  /* TG68KdotC_Kernel.vhd:1787:49  */
  assign n2529 = n2506 ? n2525 : n2501;
  /* TG68KdotC_Kernel.vhd:1787:49  */
  assign n2531 = n2506 ? n2527 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1795:58  */
  assign n2532 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1795:71  */
  assign n2534 = n2532 == 3'b010;
  /* TG68KdotC_Kernel.vhd:1795:87  */
  assign n2535 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1795:100  */
  assign n2537 = n2535 == 3'b011;
  /* TG68KdotC_Kernel.vhd:1795:78  */
  assign n2538 = n2534 | n2537;
  /* TG68KdotC_Kernel.vhd:1796:66  */
  assign n2539 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1796:78  */
  assign n2541 = n2539 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1796:95  */
  assign n2542 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1796:107  */
  assign n2544 = n2542 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1796:86  */
  assign n2545 = n2541 | n2544;
  /* TG68KdotC_Kernel.vhd:1796:57  */
  assign n2548 = n2545 ? n2528 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1796:57  */
  assign n2550 = n2545 ? n2529 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1796:57  */
  assign n2552 = n2545 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1795:49  */
  assign n2553 = n2538 ? n2548 : n2528;
  /* TG68KdotC_Kernel.vhd:1795:49  */
  assign n2554 = n2538 ? n2550 : n2529;
  /* TG68KdotC_Kernel.vhd:1795:49  */
  assign n2556 = n2538 ? n2552 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1803:58  */
  assign n2557 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1803:71  */
  assign n2559 = n2557 == 3'b101;
  /* TG68KdotC_Kernel.vhd:1804:66  */
  assign n2560 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1804:78  */
  assign n2562 = n2560 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1804:95  */
  assign n2563 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:1804:107  */
  assign n2565 = n2563 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1804:86  */
  assign n2566 = n2562 | n2565;
  /* TG68KdotC_Kernel.vhd:1804:123  */
  assign n2567 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:1804:135  */
  assign n2569 = n2567 == 3'b100;
  /* TG68KdotC_Kernel.vhd:1804:152  */
  assign n2570 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1804:155  */
  assign n2571 = ~n2570;
  /* TG68KdotC_Kernel.vhd:1804:142  */
  assign n2572 = n2571 & n2569;
  /* TG68KdotC_Kernel.vhd:1804:113  */
  assign n2573 = n2566 | n2572;
  /* TG68KdotC_Kernel.vhd:1804:57  */
  assign n2576 = n2573 ? n2553 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1804:57  */
  assign n2578 = n2573 ? n2554 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1804:57  */
  assign n2580 = n2573 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1803:49  */
  assign n2581 = n2559 ? n2576 : n2553;
  /* TG68KdotC_Kernel.vhd:1803:49  */
  assign n2582 = n2559 ? n2578 : n2554;
  /* TG68KdotC_Kernel.vhd:1803:49  */
  assign n2584 = n2559 ? n2580 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1811:58  */
  assign n2585 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1811:71  */
  assign n2587 = n2585 == 3'b110;
  /* TG68KdotC_Kernel.vhd:1812:66  */
  assign n2588 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1812:78  */
  assign n2590 = n2588 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1812:95  */
  assign n2591 = opcode[2]; // extract
  /* TG68KdotC_Kernel.vhd:1812:98  */
  assign n2592 = ~n2591;
  /* TG68KdotC_Kernel.vhd:1812:86  */
  assign n2593 = n2590 | n2592;
  /* TG68KdotC_Kernel.vhd:1812:57  */
  assign n2596 = n2593 ? n2581 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1812:57  */
  assign n2598 = n2593 ? n2582 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1812:57  */
  assign n2600 = n2593 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1811:49  */
  assign n2601 = n2587 ? n2596 : n2581;
  /* TG68KdotC_Kernel.vhd:1811:49  */
  assign n2602 = n2587 ? n2598 : n2582;
  /* TG68KdotC_Kernel.vhd:1811:49  */
  assign n2604 = n2587 ? n2600 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1819:61  */
  assign n2605 = set_exec[5]; // extract
  /* TG68KdotC_Kernel.vhd:1819:80  */
  assign n2606 = set_exec[6]; // extract
  /* TG68KdotC_Kernel.vhd:1819:69  */
  assign n2607 = n2605 | n2606;
  /* TG68KdotC_Kernel.vhd:1819:100  */
  assign n2608 = set_exec[3]; // extract
  /* TG68KdotC_Kernel.vhd:1819:89  */
  assign n2609 = n2607 | n2608;
  /* TG68KdotC_Kernel.vhd:1819:120  */
  assign n2610 = set_exec[7]; // extract
  /* TG68KdotC_Kernel.vhd:1819:109  */
  assign n2611 = n2609 | n2610;
  /* TG68KdotC_Kernel.vhd:1819:140  */
  assign n2612 = set_exec[8]; // extract
  /* TG68KdotC_Kernel.vhd:1819:129  */
  assign n2613 = n2611 | n2612;
  /* TG68KdotC_Kernel.vhd:1820:66  */
  assign n2614 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1820:69  */
  assign n2615 = ~n2614;
  /* TG68KdotC_Kernel.vhd:1820:84  */
  assign n2616 = opcode[5:0]; // extract
  /* TG68KdotC_Kernel.vhd:1820:96  */
  assign n2618 = n2616 == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1820:74  */
  assign n2619 = n2618 & n2615;
  /* TG68KdotC_Kernel.vhd:1820:119  */
  assign n2620 = set_exec[6]; // extract
  /* TG68KdotC_Kernel.vhd:1820:139  */
  assign n2621 = set_exec[5]; // extract
  /* TG68KdotC_Kernel.vhd:1820:128  */
  assign n2622 = n2620 | n2621;
  /* TG68KdotC_Kernel.vhd:1820:158  */
  assign n2623 = set_exec[7]; // extract
  /* TG68KdotC_Kernel.vhd:1820:147  */
  assign n2624 = n2622 | n2623;
  /* TG68KdotC_Kernel.vhd:1820:106  */
  assign n2625 = n2624 & n2619;
  /* TG68KdotC_Kernel.vhd:1821:92  */
  assign n2626 = ~svmode;
  /* TG68KdotC_Kernel.vhd:1821:82  */
  assign n2627 = n2626 & decodeopc;
  /* TG68KdotC_Kernel.vhd:1821:107  */
  assign n2628 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:1821:97  */
  assign n2629 = n2628 & n2627;
  /* TG68KdotC_Kernel.vhd:1827:90  */
  assign n2631 = opcode[6]; // extract
  assign n2633 = n1788[52]; // extract
  /* TG68KdotC_Kernel.vhd:1827:81  */
  assign n2634 = n2631 ? 1'b1 : n2633;
  /* TG68KdotC_Kernel.vhd:1831:104  */
  assign n2636 = set_exec[6]; // extract
  /* TG68KdotC_Kernel.vhd:1832:104  */
  assign n2637 = set_exec[7]; // extract
  /* TG68KdotC_Kernel.vhd:1833:103  */
  assign n2638 = set_exec[5]; // extract
  /* TG68KdotC_Kernel.vhd:1826:73  */
  assign n2640 = decodeopc ? 2'b01 : n1903;
  assign n2641 = {n2638, n2637, n2636};
  assign n2642 = {n2634, 1'b1};
  assign n2643 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1826:73  */
  assign n2644 = decodeopc ? n2641 : n2643;
  assign n2645 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1826:73  */
  assign n2646 = decodeopc ? n2642 : n2645;
  /* TG68KdotC_Kernel.vhd:1826:73  */
  assign n2648 = decodeopc ? 7'b0011000 : n2057;
  /* TG68KdotC_Kernel.vhd:1821:65  */
  assign n2649 = n2629 ? n1903 : n2640;
  /* TG68KdotC_Kernel.vhd:1821:65  */
  assign n2652 = n2629 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1821:65  */
  assign n2654 = n2629 ? 1'b1 : n2602;
  assign n2655 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1821:65  */
  assign n2656 = n2629 ? n2655 : n2644;
  assign n2657 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1821:65  */
  assign n2658 = n2629 ? n2657 : 1'b1;
  assign n2659 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1821:65  */
  assign n2660 = n2629 ? n2659 : n2646;
  /* TG68KdotC_Kernel.vhd:1821:65  */
  assign n2661 = n2629 ? n2057 : n2648;
  /* TG68KdotC_Kernel.vhd:1838:69  */
  assign n2662 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1838:72  */
  assign n2663 = ~n2662;
  /* TG68KdotC_Kernel.vhd:1838:86  */
  assign n2664 = opcode[5:0]; // extract
  /* TG68KdotC_Kernel.vhd:1838:98  */
  assign n2666 = n2664 != 6'b111100;
  /* TG68KdotC_Kernel.vhd:1838:77  */
  assign n2667 = n2663 | n2666;
  /* TG68KdotC_Kernel.vhd:1838:121  */
  assign n2668 = set_exec[6]; // extract
  /* TG68KdotC_Kernel.vhd:1838:141  */
  assign n2669 = set_exec[5]; // extract
  /* TG68KdotC_Kernel.vhd:1838:130  */
  assign n2670 = n2668 | n2669;
  /* TG68KdotC_Kernel.vhd:1838:160  */
  assign n2671 = set_exec[7]; // extract
  /* TG68KdotC_Kernel.vhd:1838:149  */
  assign n2672 = n2670 | n2671;
  /* TG68KdotC_Kernel.vhd:1838:169  */
  assign n2673 = ~n2672;
  /* TG68KdotC_Kernel.vhd:1838:109  */
  assign n2674 = n2667 | n2673;
  /* TG68KdotC_Kernel.vhd:1844:84  */
  assign n2678 = datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2680 = n2729 ? 1'b1 : n2048;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2682 = n2718 ? 1'b1 : n2031;
  assign n2683 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2684 = n2724 ? 1'b1 : n2683;
  assign n2685 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2686 = n2728 ? 1'b1 : n2685;
  /* TG68KdotC_Kernel.vhd:1839:65  */
  assign n2687 = n2678 & decodeopc;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2689 = n2734 ? 7'b0011101 : n2057;
  /* TG68KdotC_Kernel.vhd:1848:74  */
  assign n2690 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1848:86  */
  assign n2692 = n2690 != 2'b00;
  /* TG68KdotC_Kernel.vhd:1848:65  */
  assign n2695 = n2692 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:74  */
  assign n2696 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1851:87  */
  assign n2698 = n2696 != 3'b110;
  /* TG68KdotC_Kernel.vhd:1852:82  */
  assign n2699 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1852:94  */
  assign n2701 = n2699 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1852:73  */
  assign n2704 = n2701 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:65  */
  assign n2707 = n2698 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:65  */
  assign n2709 = n2698 ? n2704 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1857:74  */
  assign n2710 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:1857:87  */
  assign n2712 = n2710 == 2'b10;
  assign n2714 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2715 = n2726 ? 1'b1 : n2714;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2717 = n2674 ? n2707 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2718 = decodeopc & n2674;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2720 = n2674 ? n2601 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2722 = n2674 ? n2602 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2724 = decodeopc & n2674;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2726 = n2712 & n2674;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2728 = decodeopc & n2674;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2729 = n2687 & n2674;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2731 = n2674 ? n2695 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2733 = n2674 ? n2709 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1838:57  */
  assign n2734 = decodeopc & n2674;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2735 = n2789 ? n2649 : n1903;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2737 = n2625 ? 1'b0 : n2717;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2738 = n2625 ? n2031 : n2682;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2739 = n2625 ? n2601 : n2720;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2741 = n2625 ? n2652 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2742 = n2625 ? n2654 : n2722;
  assign n2743 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2744 = n2800 ? n2656 : n2743;
  assign n2745 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2746 = n2625 ? n2745 : n2684;
  assign n2747 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2748 = n2804 ? n2658 : n2747;
  assign n2749 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2750 = n2806 ? n2660 : n2749;
  assign n2751 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2752 = n2625 ? n2751 : n2715;
  assign n2753 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2754 = n2625 ? n2753 : n2686;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2755 = n2625 ? n2048 : n2680;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2757 = n2625 ? 1'b0 : n2731;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2759 = n2625 ? 1'b0 : n2733;
  /* TG68KdotC_Kernel.vhd:1820:57  */
  assign n2760 = n2625 ? n2661 : n2689;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2761 = n2625 & n2613;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2763 = n2613 ? n2737 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2764 = n2792 ? n2738 : n2031;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2766 = n2613 ? n2739 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2768 = n2613 ? n2741 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2770 = n2613 ? n2742 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2772 = n2625 & n2613;
  assign n2773 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2774 = n2802 ? n2746 : n2773;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2776 = n2625 & n2613;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2778 = n2625 & n2613;
  assign n2779 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2780 = n2808 ? n2752 : n2779;
  assign n2781 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2782 = n2810 ? n2754 : n2781;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2783 = n2811 ? n2755 : n2048;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2785 = n2613 ? n2757 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1819:49  */
  assign n2787 = n2613 ? n2759 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2788 = n2821 ? n2760 : n2057;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2789 = n2761 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2791 = n2471 ? n2763 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2792 = n2613 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2794 = n2471 ? n2766 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2796 = n2471 ? n2768 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2798 = n2471 ? n2770 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2800 = n2772 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2802 = n2613 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2804 = n2776 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2806 = n2778 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2808 = n2613 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2810 = n2613 & n2471;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2811 = n2613 & n2471;
  assign n2812 = {n2604, n2584, n2531, n2503};
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2814 = n2471 ? n2556 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2816 = n2471 ? n2812 : 4'b0000;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2818 = n2471 ? n2785 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2820 = n2471 ? n2787 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:41  */
  assign n2821 = n2613 & n2471;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2822 = n2437 ? n1903 : n2735;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2824 = n2437 ? 1'b0 : n2791;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2825 = n2437 ? n2031 : n2764;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2826 = n2437 ? n2462 : n2794;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2827 = n2437 ? n2464 : n2796;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2829 = n2437 ? 1'b1 : n2798;
  assign n2830 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2831 = n2437 ? n2830 : n2744;
  assign n2832 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2833 = n2437 ? n2832 : n2774;
  assign n2834 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2835 = n2437 ? n2834 : n2748;
  assign n2836 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2837 = n2437 ? n2836 : n2750;
  assign n2838 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2839 = n2437 ? n2838 : n2780;
  assign n2840 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2841 = n2437 ? n2840 : n2782;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2842 = n2437 ? n2048 : n2783;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2844 = n2437 ? 1'b0 : n2814;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2846 = n2437 ? 4'b0000 : n2816;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2848 = n2437 ? 1'b0 : n2818;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2850 = n2437 ? 1'b0 : n2820;
  /* TG68KdotC_Kernel.vhd:1763:33  */
  assign n2851 = n2437 ? n2057 : n2788;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2852 = n2191 & n2190;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2853 = n2190 ? n2407 : n2822;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2855 = n2190 ? 1'b0 : n2824;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2857 = n2190 ? n2409 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2858 = n2190 ? n2031 : n2825;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2859 = n2190 ? n2411 : n2826;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2861 = n2190 ? 1'b0 : n2827;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2862 = n2190 ? n2413 : n2829;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2864 = n2190 ? n2415 : 1'b0;
  assign n2865 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2866 = n2190 ? n2865 : n2831;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2868 = n2419 & n2190;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2870 = n2191 & n2190;
  assign n2871 = n2423[0]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2872 = n2190 ? n2871 : n2833;
  assign n2873 = n2423[1]; // extract
  assign n2874 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2875 = n2190 ? n2873 : n2874;
  assign n2876 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2877 = n2190 ? n2876 : n2835;
  assign n2878 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2879 = n2190 ? n2878 : n2837;
  assign n2880 = n2425[0]; // extract
  assign n2881 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2882 = n2190 ? n2880 : n2881;
  assign n2883 = n2425[1]; // extract
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2884 = n2190 ? n2883 : n2839;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2885 = n2190 ? n2427 : n2841;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2886 = n2190 ? n2048 : n2842;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2888 = n2191 & n2190;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2890 = n2431 & n2190;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2892 = n2433 & n2190;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2894 = n2190 ? 1'b0 : n2844;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2896 = n2190 ? 4'b0000 : n2846;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2898 = n2190 ? 1'b0 : n2848;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2900 = n2190 ? 1'b0 : n2850;
  /* TG68KdotC_Kernel.vhd:1696:33  */
  assign n2901 = n2190 ? n2434 : n2851;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2902 = n2095 ? n2166 : n2406;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2903 = n2095 ? n1903 : n2853;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2904 = n2095 ? n2168 : n2855;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2906 = n2095 ? 1'b0 : n2857;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2907 = n2095 ? n2031 : n2858;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2908 = n2095 ? n2171 : n2859;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2910 = n2095 ? 1'b0 : n2861;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2911 = n2095 ? n2174 : n2862;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2913 = n2095 ? n2176 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2915 = n2095 ? 1'b0 : n2864;
  assign n2916 = {n2875, n2872};
  assign n2917 = {n2884, n2882};
  assign n2918 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2919 = n2095 ? n2918 : n2866;
  assign n2920 = n1788[26]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2921 = n2095 ? n2920 : n2290;
  assign n2922 = n1788[39]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2923 = n2095 ? n2922 : n2421;
  assign n2924 = n2916[0]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2925 = n2095 ? n2153 : n2924;
  assign n2926 = n2916[1]; // extract
  assign n2927 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2928 = n2095 ? n2927 : n2926;
  assign n2929 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2930 = n2095 ? n2929 : n2877;
  assign n2931 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2932 = n2095 ? n2931 : n2879;
  assign n2933 = n1788[56:55]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2934 = n2095 ? n2933 : n2917;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2935 = n2095 ? n2155 : n2885;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2936 = n2095 ? n2048 : n2886;
  assign n2937 = n1788[82]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2938 = n2095 ? n2937 : n2429;
  assign n2939 = n1788[84]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2940 = n2095 ? n2939 : n2298;
  assign n2941 = n1788[86]; // extract
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2942 = n2095 ? n2941 : n2300;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2944 = n2095 ? 1'b0 : n2894;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2946 = n2095 ? 4'b0000 : n2896;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2948 = n2095 ? n2182 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2949 = n2095 ? n2184 : n2898;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2950 = n2095 ? n2186 : n2900;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2951 = n2095 ? n2157 : n2901;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2953 = n2063 ? 2'b00 : n2902;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2954 = n2063 ? n1903 : n2903;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2956 = n2063 ? 1'b0 : n2904;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2958 = n2063 ? 1'b0 : n2906;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2960 = n2063 ? n2090 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2961 = n2063 ? n2083 : n2907;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2963 = n2063 ? 1'b0 : n2908;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2965 = n2063 ? 1'b0 : n2910;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2967 = n2063 ? 1'b0 : n2911;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2969 = n2063 ? 1'b0 : n2913;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2971 = n2063 ? 1'b0 : n2915;
  assign n2972 = {n2928, n2925};
  assign n2973 = {1'b1, 1'b1};
  assign n2974 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2975 = n2063 ? n2974 : n2919;
  assign n2976 = n1788[26]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2977 = n2063 ? n2976 : n2921;
  assign n2978 = n1788[37]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2979 = n2063 ? n2079 : n2978;
  assign n2980 = n1788[39]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2981 = n2063 ? n2980 : n2923;
  assign n2982 = n1788[43:42]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2983 = n2063 ? n2982 : n2972;
  assign n2984 = n2973[0]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2985 = n2063 ? n2984 : n2930;
  assign n2986 = n2973[1]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2987 = n2063 ? n2986 : n2045;
  assign n2988 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2989 = n2063 ? n2988 : n2932;
  assign n2990 = n1788[56:55]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2991 = n2063 ? n2990 : n2934;
  assign n2992 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2993 = n2063 ? n2992 : n2935;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2994 = n2063 ? n2048 : n2936;
  assign n2995 = n1788[82]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2996 = n2063 ? n2995 : n2938;
  assign n2997 = n1788[84]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n2998 = n2063 ? n2997 : n2940;
  assign n2999 = n1788[86]; // extract
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3000 = n2063 ? n2999 : n2942;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3002 = n2063 ? n2074 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3004 = n2063 ? 1'b0 : n2944;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3006 = n2063 ? 4'b0000 : n2946;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3008 = n2063 ? 1'b0 : n2948;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3010 = n2063 ? 1'b0 : n2949;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3011 = n2063 ? n2076 : n2950;
  /* TG68KdotC_Kernel.vhd:1643:25  */
  assign n3012 = n2063 ? n2087 : n2951;
  /* TG68KdotC_Kernel.vhd:1642:25  */
  assign n3014 = n2058 == 4'b0000;
  /* TG68KdotC_Kernel.vhd:1877:44  */
  assign n3015 = opcode[11:10]; // extract
  /* TG68KdotC_Kernel.vhd:1877:58  */
  assign n3017 = n3015 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1877:73  */
  assign n3018 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:1877:85  */
  assign n3020 = n3018 != 3'b111;
  /* TG68KdotC_Kernel.vhd:1877:64  */
  assign n3021 = n3017 | n3020;
  /* TG68KdotC_Kernel.vhd:1878:43  */
  assign n3022 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:1878:55  */
  assign n3024 = n3022 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1878:73  */
  assign n3025 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:1878:85  */
  assign n3027 = n3025 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1878:64  */
  assign n3028 = n3024 | n3027;
  /* TG68KdotC_Kernel.vhd:1877:94  */
  assign n3029 = n3028 & n3021;
  /* TG68KdotC_Kernel.vhd:1879:43  */
  assign n3030 = opcode[13]; // extract
  /* TG68KdotC_Kernel.vhd:1879:62  */
  assign n3031 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:1879:74  */
  assign n3033 = n3031 != 3'b001;
  /* TG68KdotC_Kernel.vhd:1879:92  */
  assign n3034 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1879:104  */
  assign n3036 = n3034 != 3'b001;
  /* TG68KdotC_Kernel.vhd:1879:82  */
  assign n3037 = n3036 & n3033;
  /* TG68KdotC_Kernel.vhd:1879:52  */
  assign n3038 = n3030 | n3037;
  /* TG68KdotC_Kernel.vhd:1878:92  */
  assign n3039 = n3038 & n3029;
  /* TG68KdotC_Kernel.vhd:1882:50  */
  assign n3041 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:1882:62  */
  assign n3043 = n3041 == 3'b001;
  assign n3045 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1882:41  */
  assign n3046 = n3043 ? 1'b1 : n3045;
  /* TG68KdotC_Kernel.vhd:1885:50  */
  assign n3047 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1885:62  */
  assign n3049 = n3047 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1886:58  */
  assign n3050 = opcode[8:7]; // extract
  /* TG68KdotC_Kernel.vhd:1886:70  */
  assign n3052 = n3050 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1886:49  */
  assign n3055 = n3052 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1885:41  */
  assign n3057 = n3049 ? n3055 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:52  */
  assign n3058 = opcode[13:12]; // extract
  /* TG68KdotC_Kernel.vhd:1891:49  */
  assign n3060 = n3058 == 2'b01;
  /* TG68KdotC_Kernel.vhd:1892:49  */
  assign n3062 = n3058 == 2'b10;
  assign n3063 = {n3062, n3060};
  /* TG68KdotC_Kernel.vhd:1890:41  */
  always @*
    case (n3063)
      2'b10: n3067 = 2'b10;
      2'b01: n3067 = 2'b00;
      default: n3067 = 2'b01;
    endcase
  /* TG68KdotC_Kernel.vhd:1896:50  */
  assign n3068 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:1896:41  */
  assign n3071 = n3068 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1900:66  */
  assign n3072 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1900:78  */
  assign n3074 = n3072 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1900:57  */
  assign n3075 = nextpass | n3074;
  /* TG68KdotC_Kernel.vhd:1902:58  */
  assign n3076 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:1902:70  */
  assign n3078 = n3076 != 3'b000;
  /* TG68KdotC_Kernel.vhd:1902:49  */
  assign n3081 = n3078 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1900:41  */
  assign n3083 = n3075 ? n3081 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1900:41  */
  assign n3086 = n3075 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1907:55  */
  assign n3088 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1907:89  */
  assign n3089 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1907:101  */
  assign n3091 = n3089 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1907:107  */
  assign n3092 = decodeopc & n3091;
  /* TG68KdotC_Kernel.vhd:1907:79  */
  assign n3093 = nextpass | n3092;
  /* TG68KdotC_Kernel.vhd:1907:61  */
  assign n3094 = n3093 & n3088;
  /* TG68KdotC_Kernel.vhd:1908:60  */
  assign n3095 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:1909:57  */
  assign n3098 = n3095 == 3'b000;
  /* TG68KdotC_Kernel.vhd:1909:67  */
  assign n3100 = n3095 == 3'b001;
  /* TG68KdotC_Kernel.vhd:1909:67  */
  assign n3101 = n3098 | n3100;
  /* TG68KdotC_Kernel.vhd:1912:74  */
  assign n3102 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:1914:82  */
  assign n3104 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1914:95  */
  assign n3106 = n3104 == 3'b111;
  /* TG68KdotC_Kernel.vhd:1912:65  */
  assign n3108 = n3111 ? 1'b1 : n2045;
  assign n3109 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:1912:65  */
  assign n3110 = n3102 ? 1'b1 : n3109;
  /* TG68KdotC_Kernel.vhd:1912:65  */
  assign n3111 = n3106 & n3102;
  /* TG68KdotC_Kernel.vhd:1918:74  */
  assign n3112 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:1920:82  */
  assign n3114 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1920:95  */
  assign n3116 = n3114 == 3'b111;
  /* TG68KdotC_Kernel.vhd:1918:65  */
  assign n3118 = n3121 ? 1'b1 : n3108;
  assign n3119 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:1918:65  */
  assign n3120 = n3112 ? 1'b1 : n3119;
  /* TG68KdotC_Kernel.vhd:1918:65  */
  assign n3121 = n3116 & n3112;
  /* TG68KdotC_Kernel.vhd:1926:76  */
  assign n3122 = ~nextpass;
  assign n3124 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:1926:65  */
  assign n3125 = n3122 ? 1'b1 : n3124;
  /* TG68KdotC_Kernel.vhd:1911:57  */
  assign n3127 = n3095 == 3'b010;
  /* TG68KdotC_Kernel.vhd:1911:67  */
  assign n3129 = n3095 == 3'b011;
  /* TG68KdotC_Kernel.vhd:1911:67  */
  assign n3130 = n3127 | n3129;
  /* TG68KdotC_Kernel.vhd:1911:73  */
  assign n3132 = n3095 == 3'b100;
  /* TG68KdotC_Kernel.vhd:1911:73  */
  assign n3133 = n3130 | n3132;
  /* TG68KdotC_Kernel.vhd:1929:57  */
  assign n3135 = n3095 == 3'b101;
  /* TG68KdotC_Kernel.vhd:1932:57  */
  assign n3137 = n3095 == 3'b110;
  /* TG68KdotC_Kernel.vhd:1936:76  */
  assign n3138 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1937:73  */
  assign n3140 = n3138 == 3'b000;
  /* TG68KdotC_Kernel.vhd:1939:73  */
  assign n3143 = n3138 == 3'b001;
  assign n3144 = {n3143, n3140};
  /* TG68KdotC_Kernel.vhd:1936:65  */
  always @*
    case (n3144)
      2'b10: n3145 = 1'b1;
      2'b01: n3145 = n2048;
      default: n3145 = n2048;
    endcase
  /* TG68KdotC_Kernel.vhd:1936:65  */
  always @*
    case (n3144)
      2'b10: n3148 = 7'b0000011;
      2'b01: n3148 = 7'b0000011;
      default: n3148 = n2057;
    endcase
  /* TG68KdotC_Kernel.vhd:1935:57  */
  assign n3150 = n3095 == 3'b111;
  assign n3151 = {n3150, n3137, n3135, n3133, n3101};
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3153 = n1903;
      5'b01000: n3153 = n1903;
      5'b00100: n3153 = n1903;
      5'b00010: n3153 = 2'b11;
      5'b00001: n3153 = n1903;
      default: n3153 = n1903;
    endcase
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3155 = n2028;
      5'b01000: n3155 = 1'b1;
      5'b00100: n3155 = n2028;
      5'b00010: n3155 = n2028;
      5'b00001: n3155 = n2028;
      default: n3155 = n2028;
    endcase
  assign n3156 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3157 = n3156;
      5'b01000: n3157 = n3156;
      5'b00100: n3157 = n3156;
      5'b00010: n3157 = n3125;
      5'b00001: n3157 = n3156;
      default: n3157 = n3156;
    endcase
  assign n3158 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3159 = n3158;
      5'b01000: n3159 = n3158;
      5'b00100: n3159 = n3158;
      5'b00010: n3159 = n3110;
      5'b00001: n3159 = n3158;
      default: n3159 = n3158;
    endcase
  assign n3160 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3161 = n3160;
      5'b01000: n3161 = n3160;
      5'b00100: n3161 = n3160;
      5'b00010: n3161 = n3120;
      5'b00001: n3161 = n3160;
      default: n3161 = n3160;
    endcase
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3162 = n2045;
      5'b01000: n3162 = n2045;
      5'b00100: n3162 = n2045;
      5'b00010: n3162 = n3118;
      5'b00001: n3162 = n2045;
      default: n3162 = n2045;
    endcase
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3163 = n3145;
      5'b01000: n3163 = n2048;
      5'b00100: n3163 = n2048;
      5'b00010: n3163 = n2048;
      5'b00001: n3163 = n2048;
      default: n3163 = n2048;
    endcase
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3164 = n3057;
      5'b01000: n3164 = n3057;
      5'b00100: n3164 = n3057;
      5'b00010: n3164 = n3057;
      5'b00001: n3164 = 1'b1;
      default: n3164 = n3057;
    endcase
  /* TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3151)
      5'b10000: n3168 = n3148;
      5'b01000: n3168 = 7'b0010011;
      5'b00100: n3168 = 7'b0000111;
      5'b00010: n3168 = 7'b0000001;
      5'b00001: n3168 = n2057;
      default: n3168 = n2057;
    endcase
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3169 = n3180 ? n3153 : n1903;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3170 = n3181 ? n3155 : n2028;
  assign n3171 = {n3161, n3159};
  assign n3172 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3173 = n3202 ? n3157 : n3172;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3174 = n3203 ? n3171 : n2043;
  /* TG68KdotC_Kernel.vhd:1907:41  */
  assign n3175 = n3094 ? n3162 : n2045;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3176 = n3207 ? n3163 : n2048;
  /* TG68KdotC_Kernel.vhd:1907:41  */
  assign n3177 = n3094 ? n3164 : n3057;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3178 = n3212 ? n3168 : n2057;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3179 = n3039 ? n3067 : n1800;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3180 = n3094 & n3039;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3181 = n3094 & n3039;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3183 = n3039 ? n3071 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3186 = n3039 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3188 = n3039 ? n3083 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3190 = n3039 ? n3086 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3193 = n3039 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3196 = n3039 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3199 = n3039 ? 1'b1 : 1'b0;
  assign n3200 = {n3175, n3046};
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3202 = n3094 & n3039;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3203 = n3094 & n3039;
  assign n3204 = n1788[49]; // extract
  assign n3205 = {n2045, n3204};
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3206 = n3039 ? n3200 : n3205;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3207 = n3094 & n3039;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3209 = n3039 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3211 = n3039 ? n3177 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1877:33  */
  assign n3212 = n3094 & n3039;
  /* TG68KdotC_Kernel.vhd:1876:25  */
  assign n3214 = n2058 == 4'b0001;
  /* TG68KdotC_Kernel.vhd:1876:36  */
  assign n3216 = n2058 == 4'b0010;
  /* TG68KdotC_Kernel.vhd:1876:36  */
  assign n3217 = n3214 | n3216;
  /* TG68KdotC_Kernel.vhd:1876:43  */
  assign n3219 = n2058 == 4'b0011;
  /* TG68KdotC_Kernel.vhd:1876:43  */
  assign n3220 = n3217 | n3219;
  /* TG68KdotC_Kernel.vhd:1953:42  */
  assign n3221 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:1954:50  */
  assign n3222 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:1955:58  */
  assign n3223 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:1955:71  */
  assign n3225 = n3223 == 3'b100;
  /* TG68KdotC_Kernel.vhd:1955:88  */
  assign n3226 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1955:100  */
  assign n3228 = n3226 == 3'b000;
  /* TG68KdotC_Kernel.vhd:1955:78  */
  assign n3229 = n3228 & n3225;
  /* TG68KdotC_Kernel.vhd:1956:66  */
  assign n3230 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1956:81  */
  assign n3231 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:1956:74  */
  assign n3232 = n3231 & n3230;
  /* TG68KdotC_Kernel.vhd:1956:57  */
  assign n3239 = n3232 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1956:57  */
  assign n3242 = n3232 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1956:57  */
  assign n3245 = n3232 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1956:57  */
  assign n3247 = n3232 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1956:57  */
  assign n3249 = n3232 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1956:57  */
  assign n3251 = n3232 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1956:57  */
  assign n3253 = n3232 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:66  */
  assign n3254 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:1968:67  */
  assign n3255 = opcode[5]; // extract
  /* TG68KdotC_Kernel.vhd:1968:84  */
  assign n3256 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:1968:96  */
  assign n3258 = n3256 == 2'b10;
  /* TG68KdotC_Kernel.vhd:1968:75  */
  assign n3259 = n3255 | n3258;
  /* TG68KdotC_Kernel.vhd:1967:74  */
  assign n3260 = n3259 & n3254;
  /* TG68KdotC_Kernel.vhd:1969:66  */
  assign n3261 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1969:78  */
  assign n3263 = n3261 != 3'b100;
  /* TG68KdotC_Kernel.vhd:1968:103  */
  assign n3264 = n3263 & n3260;
  /* TG68KdotC_Kernel.vhd:1969:96  */
  assign n3265 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:1969:108  */
  assign n3267 = n3265 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1969:86  */
  assign n3268 = n3267 & n3264;
  /* TG68KdotC_Kernel.vhd:1976:74  */
  assign n3272 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1976:86  */
  assign n3274 = n3272 == 3'b010;
  /* TG68KdotC_Kernel.vhd:1976:65  */
  assign n3277 = n3274 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1976:65  */
  assign n3280 = n3274 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1976:65  */
  assign n3283 = n3274 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1982:71  */
  assign n3284 = set[62]; // extract
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3286 = n3293 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3288 = n3307 ? 1'b1 : n2031;
  /* TG68KdotC_Kernel.vhd:1986:65  */
  assign n3290 = setexecopc ? 1'b1 : n3277;
  /* TG68KdotC_Kernel.vhd:1986:65  */
  assign n3292 = setexecopc ? 1'b1 : n3280;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3293 = n3284 & n3268;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3296 = n3268 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3299 = n3268 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3302 = n3268 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3304 = n3268 ? n3290 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3306 = n3268 ? n3292 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3307 = n3284 & n3268;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3310 = n3268 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3313 = n3268 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3315 = n3268 ? n3283 : 1'b0;
  assign n3316 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3317 = n3268 ? 1'b1 : n3316;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3319 = n3268 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:57  */
  assign n3321 = n3268 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3322 = n3229 ? n1903 : n3286;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3324 = n3229 ? 1'b0 : n3296;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3326 = n3229 ? 1'b0 : n3299;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3327 = n3229 ? n3239 : n3302;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3329 = n3229 ? 1'b0 : n3304;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3331 = n3229 ? 1'b0 : n3306;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3332 = n3229 ? n2031 : n3288;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3333 = n3229 ? n3242 : n3310;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3334 = n3229 ? n3245 : n3313;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3336 = n3229 ? 1'b0 : n3315;
  assign n3337 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3338 = n3229 ? n3337 : n3317;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3339 = n3229 ? n3247 : n3319;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3341 = n3229 ? n3249 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3342 = n3229 ? n3251 : n3321;
  /* TG68KdotC_Kernel.vhd:1955:49  */
  assign n3344 = n3229 ? n3253 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1996:58  */
  assign n3345 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:1996:70  */
  assign n3347 = n3345 != 3'b001;
  /* TG68KdotC_Kernel.vhd:1997:59  */
  assign n3348 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:1997:71  */
  assign n3350 = n3348 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1997:89  */
  assign n3351 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:1997:101  */
  assign n3353 = n3351 == 2'b00;
  /* TG68KdotC_Kernel.vhd:1997:80  */
  assign n3354 = n3350 | n3353;
  /* TG68KdotC_Kernel.vhd:1996:78  */
  assign n3355 = n3354 & n3347;
  /* TG68KdotC_Kernel.vhd:1998:66  */
  assign n3356 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:2001:74  */
  assign n3358 = c_out[1]; // extract
  /* TG68KdotC_Kernel.vhd:2001:77  */
  assign n3359 = ~n3358;
  /* TG68KdotC_Kernel.vhd:2001:91  */
  assign n3360 = op1out[15]; // extract
  /* TG68KdotC_Kernel.vhd:2001:82  */
  assign n3361 = n3359 | n3360;
  /* TG68KdotC_Kernel.vhd:2001:109  */
  assign n3362 = op2out[15]; // extract
  /* TG68KdotC_Kernel.vhd:2001:100  */
  assign n3363 = n3361 | n3362;
  /* TG68KdotC_Kernel.vhd:2001:127  */
  assign n3364 = exec[31]; // extract
  /* TG68KdotC_Kernel.vhd:2001:119  */
  assign n3365 = n3364 & n3363;
  /* TG68KdotC_Kernel.vhd:2001:65  */
  assign n3368 = n3365 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2004:66  */
  assign n3369 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:2007:74  */
  assign n3371 = c_out[2]; // extract
  /* TG68KdotC_Kernel.vhd:2007:77  */
  assign n3372 = ~n3371;
  /* TG68KdotC_Kernel.vhd:2007:91  */
  assign n3373 = op1out[31]; // extract
  /* TG68KdotC_Kernel.vhd:2007:82  */
  assign n3374 = n3372 | n3373;
  /* TG68KdotC_Kernel.vhd:2007:109  */
  assign n3375 = op2out[31]; // extract
  /* TG68KdotC_Kernel.vhd:2007:100  */
  assign n3376 = n3374 | n3375;
  /* TG68KdotC_Kernel.vhd:2007:127  */
  assign n3377 = exec[31]; // extract
  /* TG68KdotC_Kernel.vhd:2007:119  */
  assign n3378 = n3377 & n3376;
  /* TG68KdotC_Kernel.vhd:2007:65  */
  assign n3381 = n3378 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2004:57  */
  assign n3383 = n3369 ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2004:57  */
  assign n3386 = n3369 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2004:57  */
  assign n3388 = n3369 ? n3381 : 1'b1;
  assign n3389 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:2004:57  */
  assign n3390 = n3369 ? 1'b1 : n3389;
  /* TG68KdotC_Kernel.vhd:1998:57  */
  assign n3392 = n3356 ? 2'b01 : n3383;
  /* TG68KdotC_Kernel.vhd:1998:57  */
  assign n3394 = n3356 ? 1'b0 : n3386;
  /* TG68KdotC_Kernel.vhd:1998:57  */
  assign n3395 = n3356 ? n3368 : n3388;
  /* TG68KdotC_Kernel.vhd:1998:57  */
  assign n3396 = n3356 ? 1'b1 : n3390;
  /* TG68KdotC_Kernel.vhd:2014:66  */
  assign n3397 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:2014:80  */
  assign n3398 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:2014:74  */
  assign n3399 = n3397 | n3398;
  /* TG68KdotC_Kernel.vhd:2015:91  */
  assign n3400 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2015:103  */
  assign n3402 = n3400 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2015:82  */
  assign n3403 = nextpass | n3402;
  /* TG68KdotC_Kernel.vhd:2015:118  */
  assign n3404 = exec[31]; // extract
  /* TG68KdotC_Kernel.vhd:2015:126  */
  assign n3405 = ~n3404;
  /* TG68KdotC_Kernel.vhd:2015:110  */
  assign n3406 = n3405 & n3403;
  /* TG68KdotC_Kernel.vhd:2015:146  */
  assign n3408 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2015:131  */
  assign n3409 = n3408 & n3406;
  /* TG68KdotC_Kernel.vhd:2015:65  */
  assign n3412 = n3409 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2020:65  */
  assign n3416 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2020:65  */
  assign n3419 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2014:57  */
  assign n3421 = n3399 ? n3416 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2014:57  */
  assign n3423 = n3399 ? n3419 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2014:57  */
  assign n3426 = n3399 ? 1'b1 : 1'b0;
  assign n3427 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3428 = n3445 ? 1'b1 : n3427;
  /* TG68KdotC_Kernel.vhd:2014:57  */
  assign n3430 = n3399 ? n3412 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3431 = n3355 ? n3392 : n1800;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3433 = n3355 ? n3421 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3435 = n3355 ? n3423 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3437 = n3355 ? n3394 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3439 = n3355 ? n3395 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3441 = n3355 ? n3426 : 1'b0;
  assign n3442 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3443 = n3355 ? n3396 : n3442;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3445 = n3399 & n3355;
  /* TG68KdotC_Kernel.vhd:1996:49  */
  assign n3447 = n3355 ? n3430 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3448 = n3222 ? n1800 : n3431;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3449 = n3222 ? n3322 : n1903;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3451 = n3222 ? n3324 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3453 = n3222 ? n3326 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3454 = n3222 ? n3327 : n3433;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3456 = n3222 ? n3329 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3457 = n3222 ? n3331 : n3435;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3458 = n3222 ? n3332 : n2031;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3459 = n3222 ? n3333 : n3437;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3460 = n3222 ? n3334 : n3439;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3461 = n3222 ? n3336 : n3441;
  assign n3462 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3463 = n3222 ? n3462 : n3443;
  assign n3464 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3465 = n3222 ? n3338 : n3464;
  assign n3466 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3467 = n3222 ? n3466 : n3428;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3469 = n3222 ? n3339 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3471 = n3222 ? n3341 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3473 = n3222 ? 1'b0 : n3447;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3475 = n3222 ? n3342 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1954:41  */
  assign n3477 = n3222 ? n3344 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2031:52  */
  assign n3478 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:2033:67  */
  assign n3479 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2033:79  */
  assign n3481 = n3479 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2034:67  */
  assign n3482 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2034:79  */
  assign n3484 = n3482 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2034:96  */
  assign n3485 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2034:108  */
  assign n3487 = n3485 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2034:87  */
  assign n3488 = n3484 | n3487;
  /* TG68KdotC_Kernel.vhd:2033:87  */
  assign n3489 = n3488 & n3481;
  /* TG68KdotC_Kernel.vhd:2035:74  */
  assign n3490 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2035:86  */
  assign n3492 = n3490 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2036:93  */
  assign n3493 = CPU[0]; // extract
  /* TG68KdotC_Kernel.vhd:2036:96  */
  assign n3494 = ~n3493;
  /* TG68KdotC_Kernel.vhd:2036:101  */
  assign n3496 = 1'b1 & n3494;
  /* TG68KdotC_Kernel.vhd:2036:86  */
  assign n3498 = 1'b0 | n3496;
  /* TG68KdotC_Kernel.vhd:2036:116  */
  assign n3499 = n3498 | svmode;
  /* TG68KdotC_Kernel.vhd:2041:87  */
  assign n3501 = CPU[0]; // extract
  /* TG68KdotC_Kernel.vhd:2041:104  */
  assign n3503 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2041:95  */
  assign n3504 = n3503 & n3501;
  /* TG68KdotC_Kernel.vhd:2041:123  */
  assign n3505 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2041:110  */
  assign n3506 = n3505 & n3504;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3508 = n3570 ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2044:90  */
  assign n3509 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2044:102  */
  assign n3511 = n3509 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2044:81  */
  assign n3514 = n3511 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2036:73  */
  assign n3515 = n3506 & n3499;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3517 = n3571 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2036:73  */
  assign n3520 = n3499 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2036:73  */
  assign n3523 = n3499 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2036:73  */
  assign n3526 = n3499 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2036:73  */
  assign n3529 = n3499 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2036:73  */
  assign n3531 = n3499 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2036:73  */
  assign n3533 = n3499 ? n3514 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2058:82  */
  assign n3537 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2058:94  */
  assign n3539 = n3537 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2058:73  */
  assign n3542 = n3539 ? 1'b1 : 1'b0;
  assign n3544 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2061:73  */
  assign n3545 = setexecopc ? 1'b1 : n3544;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3546 = n3515 & n3492;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3547 = n3499 & n3492;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3549 = n3492 ? n3520 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3552 = n3492 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3554 = n3492 ? n3523 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3556 = n3492 ? n3526 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3558 = n3492 ? n3529 : 1'b1;
  assign n3559 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3560 = n3492 ? n3559 : n3545;
  assign n3561 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3562 = n3492 ? n3561 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3564 = n3492 ? n3531 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3566 = n3492 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3568 = n3492 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2035:65  */
  assign n3569 = n3492 ? n3533 : n3542;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3570 = n3546 & n3489;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3571 = n3547 & n3489;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3573 = n3489 ? n3549 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3575 = n3489 ? n3552 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3578 = n3489 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3580 = n3489 ? n3554 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3582 = n3489 ? n3556 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3584 = n3489 ? n3558 : 1'b0;
  assign n3585 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3586 = n3489 ? n3560 : n3585;
  assign n3587 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3588 = n3489 ? n3562 : n3587;
  assign n3589 = {n3566, n3564};
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3591 = n3489 ? n3589 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3593 = n3489 ? n3568 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:57  */
  assign n3595 = n3489 ? n3569 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2032:49  */
  assign n3597 = n3478 == 3'b000;
  /* TG68KdotC_Kernel.vhd:2070:67  */
  assign n3598 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2070:79  */
  assign n3600 = n3598 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2071:67  */
  assign n3601 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2071:79  */
  assign n3603 = n3601 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2071:96  */
  assign n3604 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2071:108  */
  assign n3606 = n3604 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2071:87  */
  assign n3607 = n3603 | n3606;
  /* TG68KdotC_Kernel.vhd:2070:87  */
  assign n3608 = n3607 & n3600;
  /* TG68KdotC_Kernel.vhd:2072:74  */
  assign n3609 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2072:86  */
  assign n3611 = n3609 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2073:93  */
  assign n3612 = CPU[0]; // extract
  /* TG68KdotC_Kernel.vhd:2073:101  */
  assign n3614 = 1'b1 & n3612;
  /* TG68KdotC_Kernel.vhd:2073:86  */
  assign n3616 = 1'b0 | n3614;
  /* TG68KdotC_Kernel.vhd:2081:90  */
  assign n3618 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2081:102  */
  assign n3620 = n3618 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2081:81  */
  assign n3623 = n3620 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3625 = n3678 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2073:73  */
  assign n3628 = n3616 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2073:73  */
  assign n3631 = n3616 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2073:73  */
  assign n3634 = n3616 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2073:73  */
  assign n3637 = n3616 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2073:73  */
  assign n3639 = n3616 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2073:73  */
  assign n3641 = n3616 ? n3623 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2092:71  */
  assign n3643 = CPU[0]; // extract
  /* TG68KdotC_Kernel.vhd:2092:88  */
  assign n3645 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2092:79  */
  assign n3646 = n3645 & n3643;
  /* TG68KdotC_Kernel.vhd:2092:107  */
  assign n3647 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2092:94  */
  assign n3648 = n3647 & n3646;
  /* TG68KdotC_Kernel.vhd:2092:65  */
  assign n3650 = n3648 ? 1'b1 : make_berr;
  assign n3652 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2095:73  */
  assign n3653 = setexecopc ? 1'b1 : n3652;
  /* TG68KdotC_Kernel.vhd:2098:82  */
  assign n3654 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2098:94  */
  assign n3656 = n3654 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2098:73  */
  assign n3659 = n3656 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3660 = n3611 ? make_berr : n3650;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3661 = n3616 & n3611;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3663 = n3611 ? n3628 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3665 = n3611 ? n3631 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3667 = n3611 ? n3634 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3669 = n3611 ? n3637 : 1'b1;
  assign n3670 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3671 = n3611 ? n3670 : n3653;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3673 = n3611 ? n3639 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3675 = n3611 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2072:65  */
  assign n3676 = n3611 ? n3641 : n3659;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3677 = n3608 ? n3660 : make_berr;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3678 = n3661 & n3608;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3680 = n3608 ? n3663 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3682 = n3608 ? n3665 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3684 = n3608 ? n3667 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3686 = n3608 ? n3669 : 1'b0;
  assign n3687 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3688 = n3608 ? n3671 : n3687;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3690 = n3608 ? n3673 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3692 = n3608 ? n3675 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2070:57  */
  assign n3694 = n3608 ? n3676 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2069:49  */
  assign n3696 = n3478 == 3'b001;
  /* TG68KdotC_Kernel.vhd:2107:66  */
  assign n3697 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2107:78  */
  assign n3699 = n3697 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2108:74  */
  assign n3700 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2108:86  */
  assign n3702 = n3700 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2109:75  */
  assign n3703 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2109:87  */
  assign n3705 = n3703 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2109:105  */
  assign n3706 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2109:117  */
  assign n3708 = n3706 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2109:96  */
  assign n3709 = n3705 | n3708;
  /* TG68KdotC_Kernel.vhd:2108:94  */
  assign n3710 = n3709 & n3702;
  /* TG68KdotC_Kernel.vhd:2113:101  */
  assign n3711 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2113:113  */
  assign n3713 = n3711 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2113:91  */
  assign n3714 = n3713 & decodeopc;
  /* TG68KdotC_Kernel.vhd:2113:129  */
  assign n3716 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2113:148  */
  assign n3717 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2113:135  */
  assign n3718 = n3717 & n3716;
  /* TG68KdotC_Kernel.vhd:2113:120  */
  assign n3719 = n3714 | n3718;
  /* TG68KdotC_Kernel.vhd:2113:154  */
  assign n3720 = n3719 | direct_data;
  assign n3722 = n1788[51]; // extract
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3723 = n3793 ? 1'b1 : n3722;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3725 = n3785 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2108:65  */
  assign n3728 = n3710 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2108:65  */
  assign n3731 = n3710 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2108:65  */
  assign n3734 = n3710 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2108:65  */
  assign n3737 = n3710 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2108:65  */
  assign n3739 = n3720 & n3710;
  /* TG68KdotC_Kernel.vhd:2121:75  */
  assign n3740 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2121:87  */
  assign n3742 = n3740 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2122:75  */
  assign n3743 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2122:87  */
  assign n3745 = n3743 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2122:104  */
  assign n3746 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2122:116  */
  assign n3748 = n3746 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2122:95  */
  assign n3749 = n3745 | n3748;
  /* TG68KdotC_Kernel.vhd:2121:95  */
  assign n3750 = n3749 & n3742;
  /* TG68KdotC_Kernel.vhd:2128:82  */
  assign n3753 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2128:94  */
  assign n3755 = n3753 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2128:73  */
  assign n3758 = n3755 ? 1'b1 : 1'b0;
  assign n3760 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3761 = n3778 ? 1'b1 : n3760;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3764 = n3750 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3767 = n3750 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3770 = n3750 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3773 = n3750 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3776 = n3750 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3778 = setexecopc & n3750;
  assign n3779 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3780 = n3750 ? 1'b1 : n3779;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3782 = n3750 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3784 = n3750 ? n3758 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3785 = n3710 & n3699;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3787 = n3699 ? 1'b0 : n3764;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3788 = n3699 ? n3728 : n3767;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3789 = n3699 ? n3731 : n3770;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3790 = n3699 ? n3734 : n3773;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3791 = n3699 ? n3737 : n3776;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3793 = n3739 & n3699;
  assign n3794 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3795 = n3699 ? n3794 : n3761;
  assign n3796 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3797 = n3699 ? n3796 : n3780;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3799 = n3699 ? 1'b0 : n3782;
  /* TG68KdotC_Kernel.vhd:2107:57  */
  assign n3801 = n3699 ? 1'b0 : n3784;
  /* TG68KdotC_Kernel.vhd:2106:49  */
  assign n3803 = n3478 == 3'b010;
  /* TG68KdotC_Kernel.vhd:2140:66  */
  assign n3804 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2140:78  */
  assign n3806 = n3804 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2141:74  */
  assign n3807 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2141:86  */
  assign n3809 = n3807 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2142:75  */
  assign n3810 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2142:87  */
  assign n3812 = n3810 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2142:105  */
  assign n3813 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2142:117  */
  assign n3815 = n3813 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2142:96  */
  assign n3816 = n3812 | n3815;
  /* TG68KdotC_Kernel.vhd:2141:94  */
  assign n3817 = n3816 & n3809;
  /* TG68KdotC_Kernel.vhd:2147:109  */
  assign n3818 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2147:121  */
  assign n3820 = n3818 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2147:99  */
  assign n3821 = n3820 & decodeopc;
  /* TG68KdotC_Kernel.vhd:2147:137  */
  assign n3823 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2147:156  */
  assign n3824 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2147:143  */
  assign n3825 = n3824 & n3823;
  /* TG68KdotC_Kernel.vhd:2147:128  */
  assign n3826 = n3821 | n3825;
  /* TG68KdotC_Kernel.vhd:2147:162  */
  assign n3827 = n3826 | direct_data;
  assign n3830 = {1'b1, 1'b1};
  assign n3831 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3832 = n3933 ? n3830 : n3831;
  /* TG68KdotC_Kernel.vhd:2151:88  */
  assign n3833 = exec[52]; // extract
  /* TG68KdotC_Kernel.vhd:2151:128  */
  assign n3834 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2151:140  */
  assign n3836 = n3834 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2151:118  */
  assign n3837 = n3836 & decodeopc;
  /* TG68KdotC_Kernel.vhd:2151:100  */
  assign n3838 = n3833 | n3837;
  /* TG68KdotC_Kernel.vhd:2151:156  */
  assign n3840 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2151:175  */
  assign n3841 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2151:162  */
  assign n3842 = n3841 & n3840;
  /* TG68KdotC_Kernel.vhd:2151:147  */
  assign n3843 = n3838 | n3842;
  /* TG68KdotC_Kernel.vhd:2151:181  */
  assign n3844 = n3843 | direct_data;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3846 = n3922 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3848 = n3921 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2143:73  */
  assign n3849 = n3844 & svmode;
  /* TG68KdotC_Kernel.vhd:2143:73  */
  assign n3852 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2143:73  */
  assign n3855 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2143:73  */
  assign n3858 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2143:73  */
  assign n3861 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2143:73  */
  assign n3863 = n3827 & svmode;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3864 = svmode & n3817;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3865 = n3849 & n3817;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3867 = n3817 ? n3852 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3870 = n3817 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3872 = n3817 ? n3855 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3874 = n3817 ? n3858 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3876 = n3817 ? n3861 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2141:65  */
  assign n3878 = n3863 & n3817;
  /* TG68KdotC_Kernel.vhd:2163:74  */
  assign n3879 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2163:86  */
  assign n3881 = n3879 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2164:75  */
  assign n3882 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2164:87  */
  assign n3884 = n3882 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2164:104  */
  assign n3885 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2164:116  */
  assign n3887 = n3885 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2164:95  */
  assign n3888 = n3884 | n3887;
  /* TG68KdotC_Kernel.vhd:2163:94  */
  assign n3889 = n3888 & n3881;
  /* TG68KdotC_Kernel.vhd:2169:82  */
  assign n3892 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2169:94  */
  assign n3894 = n3892 == 3'b000;
  /* TG68KdotC_Kernel.vhd:2169:73  */
  assign n3897 = n3894 ? 1'b1 : 1'b0;
  assign n3899 = n1788[53]; // extract
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3900 = n3914 ? 1'b1 : n3899;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3903 = n3889 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3906 = n3889 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3909 = n3889 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3912 = n3889 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3914 = setexecopc & n3889;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3916 = n3889 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3918 = n3889 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2163:65  */
  assign n3920 = n3889 ? n3897 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3921 = n3864 & n3806;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3922 = n3865 & n3806;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3924 = n3806 ? 1'b0 : n3903;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3926 = n3806 ? n3867 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3927 = n3806 ? n3870 : n3906;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3929 = n3806 ? n3872 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3930 = n3806 ? n3874 : n3909;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3931 = n3806 ? n3876 : n3912;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3933 = n3878 & n3806;
  assign n3934 = n1788[53]; // extract
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3935 = n3806 ? n3934 : n3900;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3937 = n3806 ? 1'b0 : n3916;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3939 = n3806 ? 1'b0 : n3918;
  /* TG68KdotC_Kernel.vhd:2140:57  */
  assign n3941 = n3806 ? 1'b0 : n3920;
  /* TG68KdotC_Kernel.vhd:2139:49  */
  assign n3943 = n3478 == 3'b011;
  /* TG68KdotC_Kernel.vhd:2181:66  */
  assign n3944 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:2182:74  */
  assign n3945 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2182:86  */
  assign n3947 = n3945 == 3'b000;
  /* TG68KdotC_Kernel.vhd:2182:103  */
  assign n3948 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:2182:107  */
  assign n3949 = ~n3948;
  /* TG68KdotC_Kernel.vhd:2182:93  */
  assign n3950 = n3949 & n3947;
  /* TG68KdotC_Kernel.vhd:2187:82  */
  assign n3954 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2187:85  */
  assign n3955 = ~n3954;
  /* TG68KdotC_Kernel.vhd:2187:73  */
  assign n3958 = n3955 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2187:73  */
  assign n3960 = n3955 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2193:83  */
  assign n3961 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:2193:103  */
  assign n3962 = opcode[5]; // extract
  /* TG68KdotC_Kernel.vhd:2193:120  */
  assign n3963 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:2193:132  */
  assign n3965 = n3963 == 2'b10;
  /* TG68KdotC_Kernel.vhd:2193:111  */
  assign n3966 = n3962 | n3965;
  /* TG68KdotC_Kernel.vhd:2194:83  */
  assign n3967 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2194:95  */
  assign n3969 = n3967 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2194:112  */
  assign n3970 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2194:124  */
  assign n3972 = n3970 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2194:103  */
  assign n3973 = n3969 | n3972;
  /* TG68KdotC_Kernel.vhd:2193:139  */
  assign n3974 = n3973 & n3966;
  /* TG68KdotC_Kernel.vhd:2193:92  */
  assign n3975 = n3961 | n3974;
  /* TG68KdotC_Kernel.vhd:2195:83  */
  assign n3976 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:2195:87  */
  assign n3977 = ~n3976;
  /* TG68KdotC_Kernel.vhd:2195:102  */
  assign n3978 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2195:114  */
  assign n3980 = n3978 != 2'b00;
  /* TG68KdotC_Kernel.vhd:2196:82  */
  assign n3981 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2196:94  */
  assign n3983 = n3981 != 3'b100;
  /* TG68KdotC_Kernel.vhd:2195:121  */
  assign n3984 = n3983 & n3980;
  /* TG68KdotC_Kernel.vhd:2197:82  */
  assign n3985 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2197:94  */
  assign n3987 = n3985 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2196:102  */
  assign n3988 = n3987 & n3984;
  /* TG68KdotC_Kernel.vhd:2195:92  */
  assign n3989 = n3977 | n3988;
  /* TG68KdotC_Kernel.vhd:2194:133  */
  assign n3990 = n3989 & n3975;
  /* TG68KdotC_Kernel.vhd:2200:90  */
  assign n3992 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2200:93  */
  assign n3993 = ~n3992;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n3995 = n4083 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2203:91  */
  assign n3996 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2203:103  */
  assign n3998 = n3996 == 3'b100;
  /* TG68KdotC_Kernel.vhd:2203:119  */
  assign n3999 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2203:131  */
  assign n4001 = n3999 == 3'b011;
  /* TG68KdotC_Kernel.vhd:2203:110  */
  assign n4002 = n3998 | n4001;
  /* TG68KdotC_Kernel.vhd:2203:148  */
  assign n4004 = state == 2'b01;
  /* TG68KdotC_Kernel.vhd:2203:139  */
  assign n4005 = n4004 & n4002;
  /* TG68KdotC_Kernel.vhd:2203:81  */
  assign n4009 = n4005 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2203:81  */
  assign n4011 = n4005 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2207:90  */
  assign n4012 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2207:102  */
  assign n4014 = n4012 == 3'b100;
  /* TG68KdotC_Kernel.vhd:2207:81  */
  assign n4018 = n4014 ? 1'b1 : 1'b0;
  assign n4019 = n1788[48]; // extract
  /* TG68KdotC_Kernel.vhd:2207:81  */
  assign n4020 = n4014 ? 1'b1 : n4019;
  /* TG68KdotC_Kernel.vhd:2211:89  */
  assign n4022 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2211:108  */
  assign n4023 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2211:95  */
  assign n4024 = n4023 & n4022;
  assign n4027 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4028 = n4098 ? 1'b1 : n4027;
  assign n4029 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4030 = n4100 ? 1'b1 : n4029;
  /* TG68KdotC_Kernel.vhd:2217:98  */
  assign n4032 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2217:110  */
  assign n4034 = n4032 == 3'b010;
  /* TG68KdotC_Kernel.vhd:2217:126  */
  assign n4035 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2217:138  */
  assign n4037 = n4035 == 3'b011;
  /* TG68KdotC_Kernel.vhd:2217:117  */
  assign n4038 = n4034 | n4037;
  /* TG68KdotC_Kernel.vhd:2217:154  */
  assign n4039 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2217:166  */
  assign n4041 = n4039 == 3'b100;
  /* TG68KdotC_Kernel.vhd:2217:145  */
  assign n4042 = n4038 | n4041;
  assign n4044 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2217:89  */
  assign n4045 = n4042 ? n4044 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2217:89  */
  assign n4048 = n4042 ? 7'b0011010 : 7'b0000001;
  assign n4049 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4050 = n4104 ? n4045 : n4049;
  assign n4051 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4052 = n4111 ? 1'b1 : n4051;
  /* TG68KdotC_Kernel.vhd:2215:81  */
  assign n4053 = decodeopc ? n4048 : n2057;
  /* TG68KdotC_Kernel.vhd:2224:87  */
  assign n4054 = set[62]; // extract
  /* TG68KdotC_Kernel.vhd:2227:106  */
  assign n4056 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:2227:110  */
  assign n4057 = ~n4056;
  /* TG68KdotC_Kernel.vhd:2227:97  */
  assign n4061 = n4057 ? 2'b11 : 2'b10;
  assign n4062 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4063 = n4102 ? 1'b1 : n4062;
  /* TG68KdotC_Kernel.vhd:2225:89  */
  assign n4066 = movem_run ? n4061 : 2'b01;
  /* TG68KdotC_Kernel.vhd:2225:89  */
  assign n4068 = n4057 & movem_run;
  assign n4069 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4070 = n4107 ? 1'b1 : n4069;
  assign n4071 = n1788[69]; // extract
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4072 = n4109 ? 1'b1 : n4071;
  /* TG68KdotC_Kernel.vhd:2224:81  */
  assign n4074 = n4082 ? 7'b0011011 : n4053;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4075 = n4084 ? n4066 : n1903;
  /* TG68KdotC_Kernel.vhd:2224:81  */
  assign n4077 = n4068 & n4054;
  /* TG68KdotC_Kernel.vhd:2224:81  */
  assign n4079 = movem_run & n4054;
  /* TG68KdotC_Kernel.vhd:2224:81  */
  assign n4081 = movem_run & n4054;
  /* TG68KdotC_Kernel.vhd:2224:81  */
  assign n4082 = movem_run & n4054;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4083 = n3993 & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4084 = n4054 & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4087 = n3990 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4089 = n3990 ? n4018 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4092 = n3990 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4095 = n3990 ? 1'b0 : 1'b1;
  assign n4096 = {1'b1, n4020};
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4098 = n4024 & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4100 = n4024 & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4102 = n4077 & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4104 = decodeopc & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4105 = n3990 ? n4096 : n2054;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4107 = n4079 & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4109 = n4081 & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4111 = decodeopc & n3990;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4113 = n3990 ? n4009 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4115 = n3990 ? n4011 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2193:73  */
  assign n4116 = n3990 ? n4074 : n2057;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4117 = n3950 ? n3958 : n3995;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4118 = n3950 ? n1903 : n4075;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4120 = n3950 ? 1'b0 : n4087;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4123 = n3950 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4125 = n3950 ? 1'b0 : n4089;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4127 = n3950 ? 1'b0 : n4092;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4129 = n3950 ? 1'b0 : n4095;
  assign n4130 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4131 = n3950 ? n4130 : n4028;
  assign n4132 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4133 = n3950 ? n4132 : n4030;
  assign n4134 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4135 = n3950 ? n4134 : n4063;
  assign n4136 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4137 = n3950 ? n4136 : n4050;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4138 = n3950 ? n2054 : n4105;
  assign n4139 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4140 = n3950 ? n4139 : n4070;
  assign n4141 = n1788[69]; // extract
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4142 = n3950 ? n4141 : n4072;
  assign n4143 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4144 = n3950 ? n4143 : n4052;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4146 = n3950 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4148 = n3950 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4150 = n3950 ? 1'b0 : n4113;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4151 = n3950 ? 1'b1 : n4115;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4153 = n3950 ? n3960 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2182:65  */
  assign n4154 = n3950 ? n2057 : n4116;
  /* TG68KdotC_Kernel.vhd:2245:74  */
  assign n4155 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:2247:82  */
  assign n4156 = opcode[8:7]; // extract
  /* TG68KdotC_Kernel.vhd:2247:94  */
  assign n4158 = n4156 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2247:110  */
  assign n4159 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2247:122  */
  assign n4161 = n4159 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2247:100  */
  assign n4162 = n4161 & n4158;
  /* TG68KdotC_Kernel.vhd:2247:141  */
  assign n4163 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2247:153  */
  assign n4165 = n4163 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2247:171  */
  assign n4166 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2247:183  */
  assign n4168 = n4166 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2247:162  */
  assign n4169 = n4165 | n4168;
  /* TG68KdotC_Kernel.vhd:2247:130  */
  assign n4170 = n4169 & n4162;
  /* TG68KdotC_Kernel.vhd:2247:190  */
  assign n4172 = 1'b1 & n4170;
  /* TG68KdotC_Kernel.vhd:2248:102  */
  assign n4173 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2248:105  */
  assign n4174 = ~n4173;
  /* TG68KdotC_Kernel.vhd:2248:133  */
  assign n4175 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:2248:141  */
  assign n4177 = 1'b1 & n4175;
  /* TG68KdotC_Kernel.vhd:2248:126  */
  assign n4179 = 1'b0 | n4177;
  /* TG68KdotC_Kernel.vhd:2248:110  */
  assign n4180 = n4179 & n4174;
  /* TG68KdotC_Kernel.vhd:2248:91  */
  assign n4181 = n4180 & n4172;
  assign n4184 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2249:81  */
  assign n4185 = decodeopc ? 1'b1 : n4184;
  assign n4186 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2249:81  */
  assign n4187 = decodeopc ? 1'b1 : n4186;
  /* TG68KdotC_Kernel.vhd:2249:81  */
  assign n4189 = decodeopc ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:2254:96  */
  assign n4191 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2254:102  */
  assign n4192 = nextpass & n4191;
  /* TG68KdotC_Kernel.vhd:2254:130  */
  assign n4193 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2254:142  */
  assign n4195 = n4193 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2254:156  */
  assign n4196 = exec[42]; // extract
  /* TG68KdotC_Kernel.vhd:2254:148  */
  assign n4197 = n4196 & n4195;
  /* TG68KdotC_Kernel.vhd:2254:120  */
  assign n4198 = n4192 | n4197;
  /* TG68KdotC_Kernel.vhd:2259:98  */
  assign n4201 = sndopc[10]; // extract
  /* TG68KdotC_Kernel.vhd:2254:81  */
  assign n4203 = n4209 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2254:81  */
  assign n4205 = n4219 ? 7'b1010100 : n4189;
  /* TG68KdotC_Kernel.vhd:2254:81  */
  assign n4209 = n4201 & n4198;
  /* TG68KdotC_Kernel.vhd:2254:81  */
  assign n4212 = n4198 ? 1'b1 : 1'b0;
  assign n4213 = n1788[20]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4214 = n4603 ? 1'b1 : n4213;
  assign n4215 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4216 = n4607 ? 1'b1 : n4215;
  assign n4217 = n1788[67]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4218 = n4621 ? 1'b1 : n4217;
  /* TG68KdotC_Kernel.vhd:2254:81  */
  assign n4219 = n4201 & n4198;
  /* TG68KdotC_Kernel.vhd:2269:85  */
  assign n4220 = opcode[8:7]; // extract
  /* TG68KdotC_Kernel.vhd:2269:97  */
  assign n4222 = n4220 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2269:113  */
  assign n4223 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2269:125  */
  assign n4225 = n4223 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2269:103  */
  assign n4226 = n4225 & n4222;
  /* TG68KdotC_Kernel.vhd:2269:144  */
  assign n4227 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2269:156  */
  assign n4229 = n4227 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2269:174  */
  assign n4230 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2269:186  */
  assign n4232 = n4230 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2269:165  */
  assign n4233 = n4229 | n4232;
  /* TG68KdotC_Kernel.vhd:2269:133  */
  assign n4234 = n4233 & n4226;
  /* TG68KdotC_Kernel.vhd:2270:84  */
  assign n4235 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2270:115  */
  assign n4236 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:2270:123  */
  assign n4238 = 1'b1 & n4236;
  /* TG68KdotC_Kernel.vhd:2270:108  */
  assign n4240 = 1'b0 | n4238;
  /* TG68KdotC_Kernel.vhd:2270:92  */
  assign n4241 = n4240 & n4235;
  /* TG68KdotC_Kernel.vhd:2271:83  */
  assign n4242 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2271:86  */
  assign n4243 = ~n4242;
  /* TG68KdotC_Kernel.vhd:2271:114  */
  assign n4244 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:2271:122  */
  assign n4246 = 1'b1 & n4244;
  /* TG68KdotC_Kernel.vhd:2271:107  */
  assign n4248 = 1'b0 | n4246;
  /* TG68KdotC_Kernel.vhd:2271:91  */
  assign n4249 = n4248 & n4243;
  /* TG68KdotC_Kernel.vhd:2270:141  */
  assign n4250 = n4241 | n4249;
  /* TG68KdotC_Kernel.vhd:2269:193  */
  assign n4251 = n4250 & n4234;
  assign n4254 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4255 = n4316 ? 1'b1 : n4254;
  assign n4256 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4257 = n4318 ? 1'b1 : n4256;
  /* TG68KdotC_Kernel.vhd:2272:81  */
  assign n4259 = decodeopc ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:2277:96  */
  assign n4261 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2277:102  */
  assign n4262 = nextpass & n4261;
  /* TG68KdotC_Kernel.vhd:2277:130  */
  assign n4263 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2277:142  */
  assign n4265 = n4263 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2277:156  */
  assign n4266 = exec[42]; // extract
  /* TG68KdotC_Kernel.vhd:2277:148  */
  assign n4267 = n4266 & n4265;
  /* TG68KdotC_Kernel.vhd:2277:120  */
  assign n4268 = n4262 | n4267;
  /* TG68KdotC_Kernel.vhd:2281:98  */
  assign n4269 = opcode[6]; // extract
  assign n4271 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2281:89  */
  assign n4272 = n4269 ? n4271 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2281:89  */
  assign n4275 = n4269 ? 7'b1010101 : 7'b1010001;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4277 = n4297 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2277:81  */
  assign n4280 = n4268 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2277:81  */
  assign n4283 = n4268 ? 1'b1 : 1'b0;
  assign n4284 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4285 = n4314 ? n4272 : n4284;
  /* TG68KdotC_Kernel.vhd:2277:81  */
  assign n4286 = n4268 ? n4275 : n4259;
  /* TG68KdotC_Kernel.vhd:2289:107  */
  assign n4287 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2289:119  */
  assign n4289 = n4287 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2289:125  */
  assign n4290 = decodeopc & n4289;
  /* TG68KdotC_Kernel.vhd:2289:97  */
  assign n4291 = nextpass | n4290;
  /* TG68KdotC_Kernel.vhd:2289:81  */
  assign n4294 = n4291 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4296 = n4251 ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4297 = n4268 & n4251;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4300 = n4251 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4302 = n4251 ? n4280 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4304 = n4251 ? n4283 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4306 = n4251 ? n4294 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4309 = n4251 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4312 = n4251 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4314 = n4268 & n4251;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4316 = decodeopc & n4251;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4318 = decodeopc & n4251;
  /* TG68KdotC_Kernel.vhd:2269:73  */
  assign n4319 = n4251 ? n4286 : n2057;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4321 = n4181 ? 2'b10 : n4296;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4322 = n4181 ? n4203 : n4277;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4324 = n4181 ? 1'b1 : n4300;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4326 = n4181 ? 1'b0 : n4302;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4327 = n4181 ? n4212 : n4304;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4329 = n4181 ? 1'b0 : n4306;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4331 = n4181 ? 1'b0 : n4309;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4333 = n4181 ? 1'b0 : n4312;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4335 = n4198 & n4181;
  assign n4336 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4337 = n4181 ? n4336 : n4285;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4339 = n4198 & n4181;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4340 = n4181 ? n4185 : n4255;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4342 = n4198 & n4181;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4343 = n4181 ? n4187 : n4257;
  /* TG68KdotC_Kernel.vhd:2247:73  */
  assign n4344 = n4181 ? n4205 : n4319;
  /* TG68KdotC_Kernel.vhd:2299:82  */
  assign n4345 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2301:90  */
  assign n4346 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2301:102  */
  assign n4348 = n4346 == 3'b000;
  /* TG68KdotC_Kernel.vhd:2304:93  */
  assign n4351 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2304:105  */
  assign n4353 = n4351 == 3'b001;
  /* TG68KdotC_Kernel.vhd:2308:99  */
  assign n4354 = opcode[5]; // extract
  /* TG68KdotC_Kernel.vhd:2308:116  */
  assign n4355 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:2308:128  */
  assign n4357 = n4355 == 2'b10;
  /* TG68KdotC_Kernel.vhd:2308:107  */
  assign n4358 = n4354 | n4357;
  /* TG68KdotC_Kernel.vhd:2309:98  */
  assign n4359 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2309:110  */
  assign n4361 = n4359 != 3'b100;
  /* TG68KdotC_Kernel.vhd:2308:135  */
  assign n4362 = n4361 & n4358;
  /* TG68KdotC_Kernel.vhd:2310:98  */
  assign n4363 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2310:110  */
  assign n4365 = n4363 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2309:118  */
  assign n4366 = n4365 & n4362;
  /* TG68KdotC_Kernel.vhd:2313:128  */
  assign n4368 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2313:113  */
  assign n4369 = n4368 & nextpass;
  /* TG68KdotC_Kernel.vhd:2313:97  */
  assign n4372 = n4369 ? 2'b11 : n1903;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4374 = n4383 ? 1'b1 : n1892;
  assign n4375 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4376 = n4397 ? 1'b1 : n4375;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4378 = n4398 ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:2319:103  */
  assign n4379 = set[62]; // extract
  /* TG68KdotC_Kernel.vhd:2319:97  */
  assign n4381 = n4379 ? 2'b01 : n4372;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4382 = n4366 ? n4381 : n1903;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4383 = n4369 & n4366;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4386 = n4366 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4389 = n4366 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4392 = n4366 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4395 = n4366 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4397 = n4369 & n4366;
  /* TG68KdotC_Kernel.vhd:2308:89  */
  assign n4398 = n4369 & n4366;
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4399 = n4353 ? n1903 : n4382;
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4400 = n4353 ? n1892 : n4374;
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4402 = n4353 ? 1'b0 : n4386;
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4404 = n4353 ? 1'b1 : n4389;
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4406 = n4353 ? 1'b1 : n4392;
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4408 = n4353 ? 1'b0 : n4395;
  assign n4409 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4410 = n4353 ? n4409 : n4376;
  /* TG68KdotC_Kernel.vhd:2304:81  */
  assign n4411 = n4353 ? n2057 : n4378;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4412 = n4348 ? n1903 : n4399;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4413 = n4348 ? n1892 : n4400;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4415 = n4348 ? 1'b0 : n4402;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4417 = n4348 ? 1'b0 : n4404;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4419 = n4348 ? 1'b0 : n4406;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4421 = n4348 ? 1'b0 : n4408;
  assign n4422 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4423 = n4348 ? n4422 : n4410;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4425 = n4348 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4427 = n4348 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2301:81  */
  assign n4428 = n4348 ? n2057 : n4411;
  /* TG68KdotC_Kernel.vhd:2328:90  */
  assign n4429 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2328:102  */
  assign n4431 = n4429 == 3'b001;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4441 = n4514 ? 1'b1 : n1892;
  /* TG68KdotC_Kernel.vhd:2333:89  */
  assign n4444 = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2333:89  */
  assign n4447 = decodeopc ? 1'b1 : 1'b0;
  assign n4448 = n1788[36]; // extract
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4449 = n4525 ? 1'b1 : n4448;
  assign n4450 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4451 = n4527 ? 1'b1 : n4450;
  assign n4452 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4453 = n4529 ? 1'b1 : n4452;
  assign n4454 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4455 = n4535 ? 1'b1 : n4454;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4456 = n4538 ? 1'b1 : n2048;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4458 = n4545 ? 7'b0100011 : n2057;
  /* TG68KdotC_Kernel.vhd:2345:98  */
  assign n4459 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2345:110  */
  assign n4461 = n4459 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2346:99  */
  assign n4462 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2346:111  */
  assign n4464 = n4462 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2346:128  */
  assign n4465 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2346:140  */
  assign n4467 = n4465 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2346:119  */
  assign n4468 = n4464 | n4467;
  /* TG68KdotC_Kernel.vhd:2345:118  */
  assign n4469 = n4468 & n4461;
  /* TG68KdotC_Kernel.vhd:2354:106  */
  assign n4474 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2354:118  */
  assign n4476 = n4474 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2354:97  */
  assign n4479 = n4476 ? 1'b1 : 1'b0;
  assign n4481 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4482 = n4499 ? 1'b1 : n4481;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4485 = n4469 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4488 = n4469 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4491 = n4469 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4494 = n4469 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4497 = n4469 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4499 = setexecopc & n4469;
  assign n4500 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4501 = n4469 ? 1'b1 : n4500;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4503 = n4469 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4505 = n4469 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4507 = n4469 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2345:89  */
  assign n4509 = n4469 ? n4479 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4511 = n4431 ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4513 = n4431 ? 1'b0 : n4485;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4514 = decodeopc & n4431;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4516 = n4431 ? n4444 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4517 = n4431 ? n4447 : n4488;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4519 = n4431 ? 1'b0 : n4491;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4521 = n4431 ? 1'b0 : n4494;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4523 = n4431 ? 1'b0 : n4497;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4525 = decodeopc & n4431;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4527 = decodeopc & n4431;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4529 = decodeopc & n4431;
  assign n4530 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4531 = n4431 ? 1'b1 : n4530;
  assign n4532 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4533 = n4431 ? n4532 : n4482;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4535 = decodeopc & n4431;
  assign n4536 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4537 = n4431 ? n4536 : n4501;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4538 = decodeopc & n4431;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4539 = n4431 ? 1'b1 : n4503;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4541 = n4431 ? 1'b0 : n4505;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4543 = n4431 ? 1'b0 : n4507;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4544 = n4431 ? 1'b1 : n4509;
  /* TG68KdotC_Kernel.vhd:2328:81  */
  assign n4545 = decodeopc & n4431;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4547 = n4345 ? 2'b10 : n4511;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4548 = n4345 ? n4412 : n1903;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4550 = n4345 ? 1'b0 : n4513;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4551 = n4345 ? n4413 : n4441;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4553 = n4345 ? n4415 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4555 = n4345 ? 1'b0 : n4516;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4557 = n4345 ? 1'b0 : n4517;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4558 = n4345 ? n4417 : n4519;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4559 = n4345 ? n4419 : n4521;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4560 = n4345 ? n4421 : n4523;
  assign n4561 = {n4537, n4455, n4533};
  assign n4562 = n1788[36]; // extract
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4563 = n4345 ? n4562 : n4449;
  assign n4564 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4565 = n4345 ? n4564 : n4451;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4566 = n4345 ? n4423 : n4453;
  assign n4567 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4568 = n4345 ? n4567 : n4531;
  assign n4569 = n1788[56:54]; // extract
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4570 = n4345 ? n4569 : n4561;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4571 = n4345 ? n2048 : n4456;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4573 = n4345 ? 1'b0 : n4539;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4575 = n4345 ? 1'b0 : n4541;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4577 = n4345 ? n4425 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4579 = n4345 ? 1'b0 : n4543;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4580 = n4345 ? n4427 : n4544;
  /* TG68KdotC_Kernel.vhd:2299:73  */
  assign n4581 = n4345 ? n4428 : n4458;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4582 = n4155 ? n4321 : n4547;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4583 = n4155 ? n4322 : n4548;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4585 = n4155 ? 1'b0 : n4550;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4586 = n4155 ? n1892 : n4551;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4588 = n4155 ? 1'b0 : n4553;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4590 = n4155 ? 1'b0 : n4555;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4591 = n4155 ? n4324 : n4557;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4593 = n4155 ? n4326 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4595 = n4155 ? n4327 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4597 = n4155 ? n4329 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4598 = n4155 ? n4331 : n4558;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4599 = n4155 ? n4333 : n4559;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4601 = n4155 ? 1'b0 : n4560;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4603 = n4335 & n4155;
  assign n4604 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4605 = n4155 ? n4337 : n4604;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4607 = n4339 & n4155;
  assign n4608 = n1788[36]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4609 = n4155 ? n4608 : n4563;
  assign n4610 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4611 = n4155 ? n4340 : n4610;
  assign n4612 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4613 = n4155 ? n4612 : n4565;
  assign n4614 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4615 = n4155 ? n4614 : n4566;
  assign n4616 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4617 = n4155 ? n4616 : n4568;
  assign n4618 = n1788[56:54]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4619 = n4155 ? n4618 : n4570;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4621 = n4342 & n4155;
  assign n4622 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4623 = n4155 ? n4343 : n4622;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4624 = n4155 ? n2048 : n4571;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4626 = n4155 ? 1'b0 : n4573;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4628 = n4155 ? 1'b0 : n4575;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4630 = n4155 ? 1'b0 : n4577;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4632 = n4155 ? 1'b0 : n4579;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4634 = n4155 ? 1'b0 : n4580;
  /* TG68KdotC_Kernel.vhd:2245:65  */
  assign n4635 = n4155 ? n4344 : n4581;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4636 = n3944 ? n4117 : n4582;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4637 = n3944 ? n4118 : n4583;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4639 = n3944 ? 1'b0 : n4585;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4640 = n3944 ? n1892 : n4586;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4641 = n3944 ? n4120 : n4588;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4643 = n3944 ? 1'b0 : n4590;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4644 = n3944 ? n4123 : n4591;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4646 = n3944 ? 1'b0 : n4593;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4648 = n3944 ? 1'b0 : n4595;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4650 = n3944 ? 1'b0 : n4597;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4652 = n3944 ? n4125 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4653 = n3944 ? n4127 : n4598;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4654 = n3944 ? n4129 : n4599;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4656 = n3944 ? 1'b0 : n4601;
  assign n4657 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4658 = n3944 ? n4131 : n4657;
  assign n4659 = n1788[20]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4660 = n3944 ? n4659 : n4214;
  assign n4661 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4662 = n3944 ? n4661 : n4605;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4663 = n3944 ? n4133 : n4216;
  assign n4664 = n1788[36]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4665 = n3944 ? n4664 : n4609;
  assign n4666 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4667 = n3944 ? n4135 : n4666;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4668 = n3944 ? n4137 : n4611;
  assign n4669 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4670 = n3944 ? n4669 : n4613;
  assign n4671 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4672 = n3944 ? n4671 : n4615;
  assign n4673 = n4138[0]; // extract
  assign n4674 = n1788[48]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4675 = n3944 ? n4673 : n4674;
  assign n4676 = n4138[1]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4677 = n3944 ? n4676 : n4617;
  assign n4678 = n4619[0]; // extract
  assign n4679 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4680 = n3944 ? n4679 : n4678;
  assign n4681 = n4619[1]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4682 = n3944 ? n4140 : n4681;
  assign n4683 = n4619[2]; // extract
  assign n4684 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4685 = n3944 ? n4684 : n4683;
  assign n4686 = n1788[67]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4687 = n3944 ? n4686 : n4218;
  assign n4688 = n1788[69]; // extract
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4689 = n3944 ? n4142 : n4688;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4690 = n3944 ? n4144 : n4623;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4691 = n3944 ? n2048 : n4624;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4693 = n3944 ? n4146 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4695 = n3944 ? 1'b0 : n4626;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4697 = n3944 ? n4148 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4699 = n3944 ? 1'b0 : n4628;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4701 = n3944 ? 1'b0 : n4630;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4703 = n3944 ? 1'b0 : n4632;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4705 = n3944 ? n4150 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4706 = n3944 ? n4151 : n4634;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4708 = n3944 ? n4153 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2181:57  */
  assign n4709 = n3944 ? n4154 : n4635;
  /* TG68KdotC_Kernel.vhd:2180:49  */
  assign n4711 = n3478 == 3'b100;
  /* TG68KdotC_Kernel.vhd:2180:59  */
  assign n4713 = n3478 == 3'b110;
  /* TG68KdotC_Kernel.vhd:2180:59  */
  assign n4714 = n4711 | n4713;
  /* TG68KdotC_Kernel.vhd:2371:66  */
  assign n4715 = opcode[7:3]; // extract
  /* TG68KdotC_Kernel.vhd:2371:78  */
  assign n4717 = n4715 == 5'b11111;
  /* TG68KdotC_Kernel.vhd:2371:97  */
  assign n4718 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2371:109  */
  assign n4720 = n4718 != 2'b00;
  /* TG68KdotC_Kernel.vhd:2371:87  */
  assign n4721 = n4720 & n4717;
  /* TG68KdotC_Kernel.vhd:2375:75  */
  assign n4722 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2375:87  */
  assign n4724 = n4722 != 2'b11;
  /* TG68KdotC_Kernel.vhd:2376:75  */
  assign n4725 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2376:87  */
  assign n4727 = n4725 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2377:75  */
  assign n4728 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2377:87  */
  assign n4730 = n4728 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2377:104  */
  assign n4731 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2377:116  */
  assign n4733 = n4731 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2377:95  */
  assign n4734 = n4730 | n4733;
  /* TG68KdotC_Kernel.vhd:2376:95  */
  assign n4735 = n4734 & n4727;
  /* TG68KdotC_Kernel.vhd:2375:94  */
  assign n4736 = n4724 | n4735;
  /* TG68KdotC_Kernel.vhd:2378:76  */
  assign n4737 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2378:88  */
  assign n4739 = n4737 != 2'b00;
  /* TG68KdotC_Kernel.vhd:2378:105  */
  assign n4740 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2378:117  */
  assign n4742 = n4740 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2378:95  */
  assign n4743 = n4739 | n4742;
  /* TG68KdotC_Kernel.vhd:2379:75  */
  assign n4744 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2379:87  */
  assign n4746 = n4744 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2379:105  */
  assign n4747 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2379:117  */
  assign n4749 = n4747 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2379:96  */
  assign n4750 = n4746 | n4749;
  /* TG68KdotC_Kernel.vhd:2378:127  */
  assign n4751 = n4750 & n4743;
  /* TG68KdotC_Kernel.vhd:2377:125  */
  assign n4752 = n4751 & n4736;
  /* TG68KdotC_Kernel.vhd:2383:90  */
  assign n4753 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:2383:81  */
  assign n4756 = n4753 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2381:73  */
  assign n4758 = setexecopc ? n4756 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2381:73  */
  assign n4761 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:82  */
  assign n4763 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2388:94  */
  assign n4765 = n4763 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2392:90  */
  assign n4766 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2392:102  */
  assign n4768 = n4766 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2392:81  */
  assign n4771 = n4768 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4773 = n4782 ? 2'b00 : n1800;
  /* TG68KdotC_Kernel.vhd:2388:73  */
  assign n4776 = n4765 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:73  */
  assign n4779 = n4765 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:73  */
  assign n4781 = n4765 ? n4771 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4782 = n4765 & n4752;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4784 = n4752 ? n4776 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4786 = n4752 ? n4779 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4788 = n4752 ? n4758 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4790 = n4752 ? n4761 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4793 = n4752 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4796 = n4752 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4799 = n4752 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4801 = n4752 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2375:65  */
  assign n4803 = n4752 ? n4781 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4804 = n4721 ? n1800 : n4773;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4806 = n4721 ? 1'b0 : n4784;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4808 = n4721 ? 1'b0 : n4786;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4810 = n4721 ? 1'b0 : n4788;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4812 = n4721 ? 1'b0 : n4790;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4814 = n4721 ? 1'b1 : n4793;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4816 = n4721 ? 1'b1 : n4796;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4818 = n4721 ? 1'b0 : n4799;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4820 = n4721 ? 1'b0 : n4801;
  /* TG68KdotC_Kernel.vhd:2371:57  */
  assign n4822 = n4721 ? 1'b0 : n4803;
  /* TG68KdotC_Kernel.vhd:2369:49  */
  assign n4824 = n3478 == 3'b101;
  /* TG68KdotC_Kernel.vhd:2420:66  */
  assign n4825 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:2421:75  */
  assign n4826 = opcode[5]; // extract
  /* TG68KdotC_Kernel.vhd:2421:92  */
  assign n4827 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:2421:104  */
  assign n4829 = n4827 == 2'b10;
  /* TG68KdotC_Kernel.vhd:2421:83  */
  assign n4830 = n4826 | n4829;
  /* TG68KdotC_Kernel.vhd:2422:74  */
  assign n4831 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2422:86  */
  assign n4833 = n4831 != 3'b100;
  /* TG68KdotC_Kernel.vhd:2421:111  */
  assign n4834 = n4833 & n4830;
  /* TG68KdotC_Kernel.vhd:2422:104  */
  assign n4835 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2422:116  */
  assign n4837 = n4835 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2422:94  */
  assign n4838 = n4837 & n4834;
  /* TG68KdotC_Kernel.vhd:2426:80  */
  assign n4839 = exec[63]; // extract
  /* TG68KdotC_Kernel.vhd:2426:73  */
  assign n4841 = n4839 ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:2429:104  */
  assign n4843 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2429:89  */
  assign n4844 = n4843 & nextpass;
  /* TG68KdotC_Kernel.vhd:2429:120  */
  assign n4845 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2429:123  */
  assign n4846 = ~n4845;
  /* TG68KdotC_Kernel.vhd:2429:110  */
  assign n4847 = n4846 & n4844;
  /* TG68KdotC_Kernel.vhd:2429:73  */
  assign n4850 = n4847 ? 2'b11 : n1903;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4852 = n4886 ? 1'b1 : n1892;
  assign n4853 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4854 = n4903 ? 1'b1 : n4853;
  /* TG68KdotC_Kernel.vhd:2429:73  */
  assign n4856 = n4847 ? 7'b0011000 : n4841;
  /* TG68KdotC_Kernel.vhd:2436:87  */
  assign n4858 = micro_state == 7'b0000101;
  /* TG68KdotC_Kernel.vhd:2436:106  */
  assign n4859 = brief[8]; // extract
  /* TG68KdotC_Kernel.vhd:2436:109  */
  assign n4860 = ~n4859;
  /* TG68KdotC_Kernel.vhd:2436:97  */
  assign n4861 = n4860 & n4858;
  /* TG68KdotC_Kernel.vhd:2436:73  */
  assign n4863 = n4861 ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2439:81  */
  assign n4865 = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:2439:73  */
  assign n4868 = n4865 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2443:79  */
  assign n4870 = set[62]; // extract
  /* TG68KdotC_Kernel.vhd:2444:88  */
  assign n4871 = exec[73]; // extract
  /* TG68KdotC_Kernel.vhd:2444:100  */
  assign n4872 = ~n4871;
  /* TG68KdotC_Kernel.vhd:2444:105  */
  assign n4873 = n4872 | long_done;
  /* TG68KdotC_Kernel.vhd:2443:73  */
  assign n4875 = n4877 ? 1'b1 : n4863;
  /* TG68KdotC_Kernel.vhd:2443:73  */
  assign n4877 = n4873 & n4870;
  /* TG68KdotC_Kernel.vhd:2443:73  */
  assign n4879 = n4870 ? 2'b01 : n4850;
  assign n4880 = n1788[63]; // extract
  /* TG68KdotC_Kernel.vhd:2443:73  */
  assign n4881 = n4870 ? 1'b1 : n4880;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4882 = n4838 ? n4875 : make_berr;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4884 = n4838 ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4885 = n4838 ? n4879 : n1903;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4886 = n4847 & n4838;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4888 = n4838 ? n4868 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4891 = n4838 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4894 = n4838 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4897 = n4838 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4900 = n4838 ? 1'b1 : 1'b0;
  assign n4901 = {1'b1, n4881};
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4903 = n4847 & n4838;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n4904 = n5426 ? n4901 : n2055;
  /* TG68KdotC_Kernel.vhd:2421:65  */
  assign n4905 = n4838 ? n4856 : n2057;
  /* TG68KdotC_Kernel.vhd:2455:76  */
  assign n4906 = opcode[6:0]; // extract
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n4908 = n4906 == 7'b1000000;
  /* TG68KdotC_Kernel.vhd:2456:87  */
  assign n4910 = n4906 == 7'b1000001;
  /* TG68KdotC_Kernel.vhd:2456:87  */
  assign n4911 = n4908 | n4910;
  /* TG68KdotC_Kernel.vhd:2456:97  */
  assign n4913 = n4906 == 7'b1000010;
  /* TG68KdotC_Kernel.vhd:2456:97  */
  assign n4914 = n4911 | n4913;
  /* TG68KdotC_Kernel.vhd:2456:107  */
  assign n4916 = n4906 == 7'b1000011;
  /* TG68KdotC_Kernel.vhd:2456:107  */
  assign n4917 = n4914 | n4916;
  /* TG68KdotC_Kernel.vhd:2456:117  */
  assign n4919 = n4906 == 7'b1000100;
  /* TG68KdotC_Kernel.vhd:2456:117  */
  assign n4920 = n4917 | n4919;
  /* TG68KdotC_Kernel.vhd:2456:127  */
  assign n4922 = n4906 == 7'b1000101;
  /* TG68KdotC_Kernel.vhd:2456:127  */
  assign n4923 = n4920 | n4922;
  /* TG68KdotC_Kernel.vhd:2456:137  */
  assign n4925 = n4906 == 7'b1000110;
  /* TG68KdotC_Kernel.vhd:2456:137  */
  assign n4926 = n4923 | n4925;
  /* TG68KdotC_Kernel.vhd:2456:147  */
  assign n4928 = n4906 == 7'b1000111;
  /* TG68KdotC_Kernel.vhd:2456:147  */
  assign n4929 = n4926 | n4928;
  /* TG68KdotC_Kernel.vhd:2456:157  */
  assign n4931 = n4906 == 7'b1001000;
  /* TG68KdotC_Kernel.vhd:2456:157  */
  assign n4932 = n4929 | n4931;
  /* TG68KdotC_Kernel.vhd:2457:87  */
  assign n4934 = n4906 == 7'b1001001;
  /* TG68KdotC_Kernel.vhd:2457:87  */
  assign n4935 = n4932 | n4934;
  /* TG68KdotC_Kernel.vhd:2457:97  */
  assign n4937 = n4906 == 7'b1001010;
  /* TG68KdotC_Kernel.vhd:2457:97  */
  assign n4938 = n4935 | n4937;
  /* TG68KdotC_Kernel.vhd:2457:107  */
  assign n4940 = n4906 == 7'b1001011;
  /* TG68KdotC_Kernel.vhd:2457:107  */
  assign n4941 = n4938 | n4940;
  /* TG68KdotC_Kernel.vhd:2457:117  */
  assign n4943 = n4906 == 7'b1001100;
  /* TG68KdotC_Kernel.vhd:2457:117  */
  assign n4944 = n4941 | n4943;
  /* TG68KdotC_Kernel.vhd:2457:127  */
  assign n4946 = n4906 == 7'b1001101;
  /* TG68KdotC_Kernel.vhd:2457:127  */
  assign n4947 = n4944 | n4946;
  /* TG68KdotC_Kernel.vhd:2457:137  */
  assign n4949 = n4906 == 7'b1001110;
  /* TG68KdotC_Kernel.vhd:2457:137  */
  assign n4950 = n4947 | n4949;
  /* TG68KdotC_Kernel.vhd:2457:147  */
  assign n4952 = n4906 == 7'b1001111;
  /* TG68KdotC_Kernel.vhd:2457:147  */
  assign n4953 = n4950 | n4952;
  /* TG68KdotC_Kernel.vhd:2466:81  */
  assign n4961 = decodeopc ? 1'b1 : n1892;
  /* TG68KdotC_Kernel.vhd:2466:81  */
  assign n4964 = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2466:81  */
  assign n4967 = decodeopc ? 1'b1 : 1'b0;
  assign n4968 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2466:81  */
  assign n4969 = decodeopc ? 1'b1 : n4968;
  assign n4970 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2466:81  */
  assign n4971 = decodeopc ? 1'b1 : n4970;
  assign n4972 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2466:81  */
  assign n4973 = decodeopc ? 1'b1 : n4972;
  /* TG68KdotC_Kernel.vhd:2466:81  */
  assign n4975 = decodeopc ? 7'b0100011 : n2057;
  /* TG68KdotC_Kernel.vhd:2461:73  */
  assign n4977 = n4906 == 7'b1010000;
  /* TG68KdotC_Kernel.vhd:2461:87  */
  assign n4979 = n4906 == 7'b1010001;
  /* TG68KdotC_Kernel.vhd:2461:87  */
  assign n4980 = n4977 | n4979;
  /* TG68KdotC_Kernel.vhd:2461:97  */
  assign n4982 = n4906 == 7'b1010010;
  /* TG68KdotC_Kernel.vhd:2461:97  */
  assign n4983 = n4980 | n4982;
  /* TG68KdotC_Kernel.vhd:2461:107  */
  assign n4985 = n4906 == 7'b1010011;
  /* TG68KdotC_Kernel.vhd:2461:107  */
  assign n4986 = n4983 | n4985;
  /* TG68KdotC_Kernel.vhd:2461:117  */
  assign n4988 = n4906 == 7'b1010100;
  /* TG68KdotC_Kernel.vhd:2461:117  */
  assign n4989 = n4986 | n4988;
  /* TG68KdotC_Kernel.vhd:2461:127  */
  assign n4991 = n4906 == 7'b1010101;
  /* TG68KdotC_Kernel.vhd:2461:127  */
  assign n4992 = n4989 | n4991;
  /* TG68KdotC_Kernel.vhd:2461:137  */
  assign n4994 = n4906 == 7'b1010110;
  /* TG68KdotC_Kernel.vhd:2461:137  */
  assign n4995 = n4992 | n4994;
  /* TG68KdotC_Kernel.vhd:2461:147  */
  assign n4997 = n4906 == 7'b1010111;
  /* TG68KdotC_Kernel.vhd:2461:147  */
  assign n4998 = n4995 | n4997;
  /* TG68KdotC_Kernel.vhd:2481:81  */
  assign n5005 = decodeopc ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2481:81  */
  assign n5007 = decodeopc ? 1'b1 : n1892;
  /* TG68KdotC_Kernel.vhd:2481:81  */
  assign n5010 = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2481:81  */
  assign n5013 = decodeopc ? 1'b1 : 1'b0;
  assign n5014 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:2481:81  */
  assign n5015 = decodeopc ? 1'b1 : n5014;
  assign n5016 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2481:81  */
  assign n5017 = decodeopc ? 1'b1 : n5016;
  /* TG68KdotC_Kernel.vhd:2481:81  */
  assign n5019 = decodeopc ? 7'b0100101 : n2057;
  /* TG68KdotC_Kernel.vhd:2476:73  */
  assign n5021 = n4906 == 7'b1011000;
  /* TG68KdotC_Kernel.vhd:2476:87  */
  assign n5023 = n4906 == 7'b1011001;
  /* TG68KdotC_Kernel.vhd:2476:87  */
  assign n5024 = n5021 | n5023;
  /* TG68KdotC_Kernel.vhd:2476:97  */
  assign n5026 = n4906 == 7'b1011010;
  /* TG68KdotC_Kernel.vhd:2476:97  */
  assign n5027 = n5024 | n5026;
  /* TG68KdotC_Kernel.vhd:2476:107  */
  assign n5029 = n4906 == 7'b1011011;
  /* TG68KdotC_Kernel.vhd:2476:107  */
  assign n5030 = n5027 | n5029;
  /* TG68KdotC_Kernel.vhd:2476:117  */
  assign n5032 = n4906 == 7'b1011100;
  /* TG68KdotC_Kernel.vhd:2476:117  */
  assign n5033 = n5030 | n5032;
  /* TG68KdotC_Kernel.vhd:2476:127  */
  assign n5035 = n4906 == 7'b1011101;
  /* TG68KdotC_Kernel.vhd:2476:127  */
  assign n5036 = n5033 | n5035;
  /* TG68KdotC_Kernel.vhd:2476:137  */
  assign n5038 = n4906 == 7'b1011110;
  /* TG68KdotC_Kernel.vhd:2476:137  */
  assign n5039 = n5036 | n5038;
  /* TG68KdotC_Kernel.vhd:2476:147  */
  assign n5041 = n4906 == 7'b1011111;
  /* TG68KdotC_Kernel.vhd:2476:147  */
  assign n5042 = n5039 | n5041;
  /* TG68KdotC_Kernel.vhd:2492:81  */
  assign n5045 = svmode ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2492:81  */
  assign n5048 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2492:81  */
  assign n5051 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2492:81  */
  assign n5054 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2492:81  */
  assign n5057 = svmode ? 1'b0 : 1'b1;
  assign n5058 = n1896[0]; // extract
  /* TG68KdotC_Kernel.vhd:2492:81  */
  assign n5059 = svmode ? 1'b1 : n5058;
  /* TG68KdotC_Kernel.vhd:2491:73  */
  assign n5061 = n4906 == 7'b1100000;
  /* TG68KdotC_Kernel.vhd:2491:87  */
  assign n5063 = n4906 == 7'b1100001;
  /* TG68KdotC_Kernel.vhd:2491:87  */
  assign n5064 = n5061 | n5063;
  /* TG68KdotC_Kernel.vhd:2491:97  */
  assign n5066 = n4906 == 7'b1100010;
  /* TG68KdotC_Kernel.vhd:2491:97  */
  assign n5067 = n5064 | n5066;
  /* TG68KdotC_Kernel.vhd:2491:107  */
  assign n5069 = n4906 == 7'b1100011;
  /* TG68KdotC_Kernel.vhd:2491:107  */
  assign n5070 = n5067 | n5069;
  /* TG68KdotC_Kernel.vhd:2491:117  */
  assign n5072 = n4906 == 7'b1100100;
  /* TG68KdotC_Kernel.vhd:2491:117  */
  assign n5073 = n5070 | n5072;
  /* TG68KdotC_Kernel.vhd:2491:127  */
  assign n5075 = n4906 == 7'b1100101;
  /* TG68KdotC_Kernel.vhd:2491:127  */
  assign n5076 = n5073 | n5075;
  /* TG68KdotC_Kernel.vhd:2491:137  */
  assign n5078 = n4906 == 7'b1100110;
  /* TG68KdotC_Kernel.vhd:2491:137  */
  assign n5079 = n5076 | n5078;
  /* TG68KdotC_Kernel.vhd:2491:147  */
  assign n5081 = n4906 == 7'b1100111;
  /* TG68KdotC_Kernel.vhd:2491:147  */
  assign n5082 = n5079 | n5081;
  /* TG68KdotC_Kernel.vhd:2504:81  */
  assign n5086 = svmode ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2504:81  */
  assign n5089 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2504:81  */
  assign n5092 = svmode ? 1'b0 : 1'b1;
  assign n5093 = n1896[1]; // extract
  /* TG68KdotC_Kernel.vhd:2504:81  */
  assign n5094 = svmode ? 1'b1 : n5093;
  /* TG68KdotC_Kernel.vhd:2504:81  */
  assign n5096 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2503:73  */
  assign n5098 = n4906 == 7'b1101000;
  /* TG68KdotC_Kernel.vhd:2503:87  */
  assign n5100 = n4906 == 7'b1101001;
  /* TG68KdotC_Kernel.vhd:2503:87  */
  assign n5101 = n5098 | n5100;
  /* TG68KdotC_Kernel.vhd:2503:97  */
  assign n5103 = n4906 == 7'b1101010;
  /* TG68KdotC_Kernel.vhd:2503:97  */
  assign n5104 = n5101 | n5103;
  /* TG68KdotC_Kernel.vhd:2503:107  */
  assign n5106 = n4906 == 7'b1101011;
  /* TG68KdotC_Kernel.vhd:2503:107  */
  assign n5107 = n5104 | n5106;
  /* TG68KdotC_Kernel.vhd:2503:117  */
  assign n5109 = n4906 == 7'b1101100;
  /* TG68KdotC_Kernel.vhd:2503:117  */
  assign n5110 = n5107 | n5109;
  /* TG68KdotC_Kernel.vhd:2503:127  */
  assign n5112 = n4906 == 7'b1101101;
  /* TG68KdotC_Kernel.vhd:2503:127  */
  assign n5113 = n5110 | n5112;
  /* TG68KdotC_Kernel.vhd:2503:137  */
  assign n5115 = n4906 == 7'b1101110;
  /* TG68KdotC_Kernel.vhd:2503:137  */
  assign n5116 = n5113 | n5115;
  /* TG68KdotC_Kernel.vhd:2503:147  */
  assign n5118 = n4906 == 7'b1101111;
  /* TG68KdotC_Kernel.vhd:2503:147  */
  assign n5119 = n5116 | n5118;
  /* TG68KdotC_Kernel.vhd:2515:90  */
  assign n5120 = ~svmode;
  /* TG68KdotC_Kernel.vhd:2520:89  */
  assign n5124 = decodeopc ? 6'b000000 : n1785;
  assign n5125 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2520:89  */
  assign n5126 = decodeopc ? 1'b1 : n5125;
  /* TG68KdotC_Kernel.vhd:2515:81  */
  assign n5127 = n5120 ? n1785 : n5124;
  /* TG68KdotC_Kernel.vhd:2515:81  */
  assign n5130 = n5120 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2515:81  */
  assign n5133 = n5120 ? 1'b1 : 1'b0;
  assign n5134 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2515:81  */
  assign n5135 = n5120 ? n5134 : n5126;
  assign n5136 = n1788[74]; // extract
  /* TG68KdotC_Kernel.vhd:2515:81  */
  assign n5137 = n5120 ? n5136 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2514:73  */
  assign n5139 = n4906 == 7'b1110000;
  /* TG68KdotC_Kernel.vhd:2526:73  */
  assign n5141 = n4906 == 7'b1110001;
  /* TG68KdotC_Kernel.vhd:2529:90  */
  assign n5142 = ~svmode;
  /* TG68KdotC_Kernel.vhd:2533:89  */
  assign n5144 = decodeopc ? 1'b1 : n2025;
  /* TG68KdotC_Kernel.vhd:2533:89  */
  assign n5147 = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2537:89  */
  assign n5149 = stop ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2529:81  */
  assign n5150 = n5142 ? make_berr : n5149;
  /* TG68KdotC_Kernel.vhd:2529:81  */
  assign n5151 = n5142 ? n2025 : n5144;
  /* TG68KdotC_Kernel.vhd:2529:81  */
  assign n5154 = n5142 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2529:81  */
  assign n5157 = n5142 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2529:81  */
  assign n5159 = n5142 ? 1'b0 : n5147;
  /* TG68KdotC_Kernel.vhd:2528:73  */
  assign n5161 = n4906 == 7'b1110010;
  /* TG68KdotC_Kernel.vhd:2544:104  */
  assign n5162 = opcode[2]; // extract
  /* TG68KdotC_Kernel.vhd:2544:95  */
  assign n5163 = svmode | n5162;
  /* TG68KdotC_Kernel.vhd:2549:106  */
  assign n5165 = opcode[2]; // extract
  assign n5168 = n1788[59]; // extract
  /* TG68KdotC_Kernel.vhd:2549:97  */
  assign n5169 = n5165 ? n5168 : 1'b1;
  assign n5170 = n1788[60]; // extract
  /* TG68KdotC_Kernel.vhd:2549:97  */
  assign n5171 = n5165 ? 1'b1 : n5170;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5173 = n5183 ? 2'b10 : n1903;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5175 = n5184 ? 1'b1 : n1892;
  assign n5176 = {n5171, n5169};
  assign n5177 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5178 = n5192 ? 1'b1 : n5177;
  assign n5179 = n1788[60:59]; // extract
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5180 = n5194 ? n5176 : n5179;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5182 = n5195 ? 7'b0101011 : n2057;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5183 = decodeopc & n5163;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5184 = decodeopc & n5163;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5187 = n5163 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5190 = n5163 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5192 = decodeopc & n5163;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5194 = decodeopc & n5163;
  /* TG68KdotC_Kernel.vhd:2544:81  */
  assign n5195 = decodeopc & n5163;
  /* TG68KdotC_Kernel.vhd:2543:73  */
  assign n5197 = n4906 == 7'b1110011;
  /* TG68KdotC_Kernel.vhd:2543:87  */
  assign n5199 = n4906 == 7'b1110111;
  /* TG68KdotC_Kernel.vhd:2543:87  */
  assign n5200 = n5197 | n5199;
  /* TG68KdotC_Kernel.vhd:2563:81  */
  assign n5205 = decodeopc ? 2'b10 : n1903;
  /* TG68KdotC_Kernel.vhd:2563:81  */
  assign n5207 = decodeopc ? 1'b1 : n1892;
  /* TG68KdotC_Kernel.vhd:2563:81  */
  assign n5209 = decodeopc ? 1'b1 : n2031;
  assign n5210 = {1'b1, 1'b1};
  assign n5211 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2563:81  */
  assign n5212 = decodeopc ? 1'b1 : n5211;
  assign n5213 = n1788[58:57]; // extract
  /* TG68KdotC_Kernel.vhd:2563:81  */
  assign n5214 = decodeopc ? n5210 : n5213;
  /* TG68KdotC_Kernel.vhd:2563:81  */
  assign n5216 = decodeopc ? 7'b0110000 : n2057;
  /* TG68KdotC_Kernel.vhd:2561:73  */
  assign n5218 = n4906 == 7'b1110100;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5223 = decodeopc ? 2'b10 : n1903;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5225 = decodeopc ? 1'b1 : n1892;
  assign n5226 = {1'b1, 1'b1};
  assign n5227 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5228 = decodeopc ? 1'b1 : n5227;
  assign n5229 = n1788[58:57]; // extract
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5230 = decodeopc ? n5226 : n5229;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5232 = decodeopc ? 7'b0011000 : n2057;
  /* TG68KdotC_Kernel.vhd:2574:73  */
  assign n5234 = n4906 == 7'b1110101;
  /* TG68KdotC_Kernel.vhd:2586:81  */
  assign n5236 = decodeopc ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2589:89  */
  assign n5237 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:2589:106  */
  assign n5239 = state == 2'b01;
  /* TG68KdotC_Kernel.vhd:2589:97  */
  assign n5240 = n5239 & n5237;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5243 = n5240 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5246 = n5240 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2585:73  */
  assign n5248 = n4906 == 7'b1110110;
  /* TG68KdotC_Kernel.vhd:2595:87  */
  assign n5250 = CPU == 2'b00;
  /* TG68KdotC_Kernel.vhd:2598:93  */
  assign n5251 = ~svmode;
  /* TG68KdotC_Kernel.vhd:2603:106  */
  assign n5252 = last_data_read[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:2603:119  */
  assign n5254 = n5252 == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:2605:106  */
  assign n5256 = opcode[0]; // extract
  assign n5258 = n1896[0]; // extract
  /* TG68KdotC_Kernel.vhd:2605:97  */
  assign n5259 = n5256 ? 1'b1 : n5258;
  assign n5260 = {1'b1, n5259};
  /* TG68KdotC_Kernel.vhd:2603:89  */
  assign n5261 = n5254 ? n5260 : n1896;
  /* TG68KdotC_Kernel.vhd:2609:98  */
  assign n5262 = opcode[0]; // extract
  /* TG68KdotC_Kernel.vhd:2609:101  */
  assign n5263 = ~n5262;
  /* TG68KdotC_Kernel.vhd:2609:89  */
  assign n5267 = n5263 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2609:89  */
  assign n5269 = n5263 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2614:89  */
  assign n5271 = decodeopc ? 1'b1 : n2028;
  /* TG68KdotC_Kernel.vhd:2614:89  */
  assign n5273 = decodeopc ? 7'b1001001 : n2057;
  /* TG68KdotC_Kernel.vhd:2598:81  */
  assign n5275 = n5251 ? n1800 : 2'b10;
  /* TG68KdotC_Kernel.vhd:2598:81  */
  assign n5276 = n5251 ? n2028 : n5271;
  /* TG68KdotC_Kernel.vhd:2598:81  */
  assign n5279 = n5251 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2598:81  */
  assign n5282 = n5251 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2598:81  */
  assign n5283 = n5251 ? n1896 : n5261;
  assign n5284 = {n5269, n5267};
  /* TG68KdotC_Kernel.vhd:2598:81  */
  assign n5286 = n5251 ? 2'b00 : n5284;
  /* TG68KdotC_Kernel.vhd:2598:81  */
  assign n5287 = n5251 ? n2057 : n5273;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5288 = n5250 ? n1800 : n5275;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5289 = n5250 ? n2028 : n5276;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5292 = n5250 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5294 = n5250 ? 1'b0 : n5279;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5296 = n5250 ? 1'b1 : n5282;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5297 = n5250 ? n1896 : n5283;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5299 = n5250 ? 2'b00 : n5286;
  /* TG68KdotC_Kernel.vhd:2595:81  */
  assign n5300 = n5250 ? n2057 : n5287;
  /* TG68KdotC_Kernel.vhd:2594:73  */
  assign n5302 = n4906 == 7'b1111010;
  /* TG68KdotC_Kernel.vhd:2594:87  */
  assign n5304 = n4906 == 7'b1111011;
  /* TG68KdotC_Kernel.vhd:2594:87  */
  assign n5305 = n5302 | n5304;
  assign n5306 = {n5305, n5248, n5234, n5218, n5200, n5161, n5141, n5139, n5119, n5082, n5042, n4998, n4953};
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5307 = make_berr;
      13'b0100000000000: n5307 = make_berr;
      13'b0010000000000: n5307 = make_berr;
      13'b0001000000000: n5307 = make_berr;
      13'b0000100000000: n5307 = make_berr;
      13'b0000010000000: n5307 = n5150;
      13'b0000001000000: n5307 = make_berr;
      13'b0000000100000: n5307 = make_berr;
      13'b0000000010000: n5307 = make_berr;
      13'b0000000001000: n5307 = make_berr;
      13'b0000000000100: n5307 = make_berr;
      13'b0000000000010: n5307 = make_berr;
      13'b0000000000001: n5307 = make_berr;
      default: n5307 = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5312 = n5288;
      13'b0100000000000: n5312 = n1800;
      13'b0010000000000: n5312 = 2'b10;
      13'b0001000000000: n5312 = 2'b10;
      13'b0000100000000: n5312 = n1800;
      13'b0000010000000: n5312 = n1800;
      13'b0000001000000: n5312 = n1800;
      13'b0000000100000: n5312 = n1800;
      13'b0000000010000: n5312 = n5086;
      13'b0000000001000: n5312 = n5045;
      13'b0000000000100: n5312 = 2'b10;
      13'b0000000000010: n5312 = 2'b10;
      13'b0000000000001: n5312 = n1800;
      default: n5312 = n1800;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5313 = n1903;
      13'b0100000000000: n5313 = n5236;
      13'b0010000000000: n5313 = n5223;
      13'b0001000000000: n5313 = n5205;
      13'b0000100000000: n5313 = n5173;
      13'b0000010000000: n5313 = n1903;
      13'b0000001000000: n5313 = n1903;
      13'b0000000100000: n5313 = n1903;
      13'b0000000010000: n5313 = n1903;
      13'b0000000001000: n5313 = n1903;
      13'b0000000000100: n5313 = n5005;
      13'b0000000000010: n5313 = n1903;
      13'b0000000000001: n5313 = n1903;
      default: n5313 = n1903;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5314 = n2025;
      13'b0100000000000: n5314 = n2025;
      13'b0010000000000: n5314 = n2025;
      13'b0001000000000: n5314 = n2025;
      13'b0000100000000: n5314 = n2025;
      13'b0000010000000: n5314 = n5151;
      13'b0000001000000: n5314 = n2025;
      13'b0000000100000: n5314 = n2025;
      13'b0000000010000: n5314 = n2025;
      13'b0000000001000: n5314 = n2025;
      13'b0000000000100: n5314 = n2025;
      13'b0000000000010: n5314 = n2025;
      13'b0000000000001: n5314 = n2025;
      default: n5314 = n2025;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5315 = n5289;
      13'b0100000000000: n5315 = n2028;
      13'b0010000000000: n5315 = n2028;
      13'b0001000000000: n5315 = n2028;
      13'b0000100000000: n5315 = n2028;
      13'b0000010000000: n5315 = n2028;
      13'b0000001000000: n5315 = n2028;
      13'b0000000100000: n5315 = n2028;
      13'b0000000010000: n5315 = n2028;
      13'b0000000001000: n5315 = n2028;
      13'b0000000000100: n5315 = n2028;
      13'b0000000000010: n5315 = n2028;
      13'b0000000000001: n5315 = n2028;
      default: n5315 = n2028;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5316 = n1892;
      13'b0100000000000: n5316 = n1892;
      13'b0010000000000: n5316 = n5225;
      13'b0001000000000: n5316 = n5207;
      13'b0000100000000: n5316 = n5175;
      13'b0000010000000: n5316 = n1892;
      13'b0000001000000: n5316 = n1892;
      13'b0000000100000: n5316 = n1892;
      13'b0000000010000: n5316 = n1892;
      13'b0000000001000: n5316 = n1892;
      13'b0000000000100: n5316 = n5007;
      13'b0000000000010: n5316 = n4961;
      13'b0000000000001: n5316 = n1892;
      default: n5316 = n1892;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5318 = 1'b0;
      13'b0100000000000: n5318 = 1'b0;
      13'b0010000000000: n5318 = 1'b0;
      13'b0001000000000: n5318 = 1'b0;
      13'b0000100000000: n5318 = 1'b0;
      13'b0000010000000: n5318 = 1'b0;
      13'b0000001000000: n5318 = 1'b0;
      13'b0000000100000: n5318 = 1'b0;
      13'b0000000010000: n5318 = 1'b0;
      13'b0000000001000: n5318 = n5048;
      13'b0000000000100: n5318 = n5010;
      13'b0000000000010: n5318 = n4964;
      13'b0000000000001: n5318 = 1'b0;
      default: n5318 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5320 = 1'b0;
      13'b0100000000000: n5320 = 1'b0;
      13'b0010000000000: n5320 = 1'b0;
      13'b0001000000000: n5320 = 1'b0;
      13'b0000100000000: n5320 = 1'b0;
      13'b0000010000000: n5320 = 1'b0;
      13'b0000001000000: n5320 = 1'b0;
      13'b0000000100000: n5320 = 1'b0;
      13'b0000000010000: n5320 = 1'b0;
      13'b0000000001000: n5320 = n5051;
      13'b0000000000100: n5320 = n5013;
      13'b0000000000010: n5320 = n4967;
      13'b0000000000001: n5320 = 1'b0;
      default: n5320 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5321 = n1785;
      13'b0100000000000: n5321 = n1785;
      13'b0010000000000: n5321 = n1785;
      13'b0001000000000: n5321 = n1785;
      13'b0000100000000: n5321 = n1785;
      13'b0000010000000: n5321 = n1785;
      13'b0000001000000: n5321 = n1785;
      13'b0000000100000: n5321 = n5127;
      13'b0000000010000: n5321 = n1785;
      13'b0000000001000: n5321 = n1785;
      13'b0000000000100: n5321 = n1785;
      13'b0000000000010: n5321 = n1785;
      13'b0000000000001: n5321 = n1785;
      default: n5321 = n1785;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5322 = n2031;
      13'b0100000000000: n5322 = n2031;
      13'b0010000000000: n5322 = n2031;
      13'b0001000000000: n5322 = n5209;
      13'b0000100000000: n5322 = n2031;
      13'b0000010000000: n5322 = n2031;
      13'b0000001000000: n5322 = n2031;
      13'b0000000100000: n5322 = n2031;
      13'b0000000010000: n5322 = n2031;
      13'b0000000001000: n5322 = n2031;
      13'b0000000000100: n5322 = n2031;
      13'b0000000000010: n5322 = n2031;
      13'b0000000000001: n5322 = n2031;
      default: n5322 = n2031;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5325 = n5292;
      13'b0100000000000: n5325 = 1'b0;
      13'b0010000000000: n5325 = 1'b0;
      13'b0001000000000: n5325 = 1'b0;
      13'b0000100000000: n5325 = 1'b0;
      13'b0000010000000: n5325 = 1'b0;
      13'b0000001000000: n5325 = 1'b0;
      13'b0000000100000: n5325 = 1'b0;
      13'b0000000010000: n5325 = 1'b0;
      13'b0000000001000: n5325 = 1'b0;
      13'b0000000000100: n5325 = 1'b0;
      13'b0000000000010: n5325 = 1'b0;
      13'b0000000000001: n5325 = 1'b0;
      default: n5325 = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5327 = n5294;
      13'b0100000000000: n5327 = 1'b0;
      13'b0010000000000: n5327 = 1'b0;
      13'b0001000000000: n5327 = 1'b0;
      13'b0000100000000: n5327 = n5187;
      13'b0000010000000: n5327 = n5154;
      13'b0000001000000: n5327 = 1'b0;
      13'b0000000100000: n5327 = n5130;
      13'b0000000010000: n5327 = n5089;
      13'b0000000001000: n5327 = n5054;
      13'b0000000000100: n5327 = 1'b0;
      13'b0000000000010: n5327 = 1'b0;
      13'b0000000000001: n5327 = 1'b0;
      default: n5327 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5330 = 1'b0;
      13'b0100000000000: n5330 = 1'b0;
      13'b0010000000000: n5330 = 1'b0;
      13'b0001000000000: n5330 = 1'b0;
      13'b0000100000000: n5330 = 1'b0;
      13'b0000010000000: n5330 = 1'b0;
      13'b0000001000000: n5330 = 1'b0;
      13'b0000000100000: n5330 = 1'b0;
      13'b0000000010000: n5330 = 1'b0;
      13'b0000000001000: n5330 = 1'b0;
      13'b0000000000100: n5330 = 1'b0;
      13'b0000000000010: n5330 = 1'b0;
      13'b0000000000001: n5330 = 1'b1;
      default: n5330 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5332 = 1'b0;
      13'b0100000000000: n5332 = n5243;
      13'b0010000000000: n5332 = 1'b0;
      13'b0001000000000: n5332 = 1'b0;
      13'b0000100000000: n5332 = 1'b0;
      13'b0000010000000: n5332 = 1'b0;
      13'b0000001000000: n5332 = 1'b0;
      13'b0000000100000: n5332 = 1'b0;
      13'b0000000010000: n5332 = 1'b0;
      13'b0000000001000: n5332 = 1'b0;
      13'b0000000000100: n5332 = 1'b0;
      13'b0000000000010: n5332 = 1'b0;
      13'b0000000000001: n5332 = 1'b0;
      default: n5332 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5336 = n5296;
      13'b0100000000000: n5336 = n5246;
      13'b0010000000000: n5336 = 1'b0;
      13'b0001000000000: n5336 = 1'b0;
      13'b0000100000000: n5336 = n5190;
      13'b0000010000000: n5336 = n5157;
      13'b0000001000000: n5336 = 1'b0;
      13'b0000000100000: n5336 = n5133;
      13'b0000000010000: n5336 = n5092;
      13'b0000000001000: n5336 = n5057;
      13'b0000000000100: n5336 = 1'b0;
      13'b0000000000010: n5336 = 1'b0;
      13'b0000000000001: n5336 = 1'b1;
      default: n5336 = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5338 = 1'b0;
      13'b0100000000000: n5338 = 1'b0;
      13'b0010000000000: n5338 = 1'b0;
      13'b0001000000000: n5338 = 1'b0;
      13'b0000100000000: n5338 = 1'b0;
      13'b0000010000000: n5338 = n5159;
      13'b0000001000000: n5338 = 1'b0;
      13'b0000000100000: n5338 = 1'b0;
      13'b0000000010000: n5338 = 1'b0;
      13'b0000000001000: n5338 = 1'b0;
      13'b0000000000100: n5338 = 1'b0;
      13'b0000000000010: n5338 = 1'b0;
      13'b0000000000001: n5338 = 1'b0;
      default: n5338 = 1'b0;
    endcase
  assign n5339 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5340 = n5339;
      13'b0100000000000: n5340 = n5339;
      13'b0010000000000: n5340 = n5339;
      13'b0001000000000: n5340 = n5339;
      13'b0000100000000: n5340 = n5339;
      13'b0000010000000: n5340 = n5339;
      13'b0000001000000: n5340 = n5339;
      13'b0000000100000: n5340 = n5339;
      13'b0000000010000: n5340 = n5339;
      13'b0000000001000: n5340 = n5339;
      13'b0000000000100: n5340 = n5015;
      13'b0000000000010: n5340 = n5339;
      13'b0000000000001: n5340 = n5339;
      default: n5340 = n5339;
    endcase
  assign n5341 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5342 = n5341;
      13'b0100000000000: n5342 = n5341;
      13'b0010000000000: n5342 = n5341;
      13'b0001000000000: n5342 = n5341;
      13'b0000100000000: n5342 = n5341;
      13'b0000010000000: n5342 = n5341;
      13'b0000001000000: n5342 = n5341;
      13'b0000000100000: n5342 = n5135;
      13'b0000000010000: n5342 = n5341;
      13'b0000000001000: n5342 = n5341;
      13'b0000000000100: n5342 = n5341;
      13'b0000000000010: n5342 = n5341;
      13'b0000000000001: n5342 = n5341;
      default: n5342 = n5341;
    endcase
  assign n5343 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5344 = n5343;
      13'b0100000000000: n5344 = n5343;
      13'b0010000000000: n5344 = n5343;
      13'b0001000000000: n5344 = n5343;
      13'b0000100000000: n5344 = n5343;
      13'b0000010000000: n5344 = n5343;
      13'b0000001000000: n5344 = n5343;
      13'b0000000100000: n5344 = n5343;
      13'b0000000010000: n5344 = n5343;
      13'b0000000001000: n5344 = n5343;
      13'b0000000000100: n5344 = n5017;
      13'b0000000000010: n5344 = n5343;
      13'b0000000000001: n5344 = n5343;
      default: n5344 = n5343;
    endcase
  assign n5345 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5346 = n5345;
      13'b0100000000000: n5346 = n5345;
      13'b0010000000000: n5346 = n5345;
      13'b0001000000000: n5346 = n5345;
      13'b0000100000000: n5346 = n5345;
      13'b0000010000000: n5346 = n5345;
      13'b0000001000000: n5346 = n5345;
      13'b0000000100000: n5346 = n5345;
      13'b0000000010000: n5346 = n5345;
      13'b0000000001000: n5346 = n5345;
      13'b0000000000100: n5346 = n5345;
      13'b0000000000010: n5346 = n4969;
      13'b0000000000001: n5346 = n5345;
      default: n5346 = n5345;
    endcase
  assign n5347 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5348 = n5347;
      13'b0100000000000: n5348 = n5347;
      13'b0010000000000: n5348 = n5228;
      13'b0001000000000: n5348 = n5212;
      13'b0000100000000: n5348 = n5178;
      13'b0000010000000: n5348 = n5347;
      13'b0000001000000: n5348 = n5347;
      13'b0000000100000: n5348 = n5347;
      13'b0000000010000: n5348 = n5347;
      13'b0000000001000: n5348 = n5347;
      13'b0000000000100: n5348 = n5347;
      13'b0000000000010: n5348 = n5347;
      13'b0000000000001: n5348 = n5347;
      default: n5348 = n5347;
    endcase
  assign n5349 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5350 = n5349;
      13'b0100000000000: n5350 = n5349;
      13'b0010000000000: n5350 = n5349;
      13'b0001000000000: n5350 = n5349;
      13'b0000100000000: n5350 = n5349;
      13'b0000010000000: n5350 = n5349;
      13'b0000001000000: n5350 = n5349;
      13'b0000000100000: n5350 = n5349;
      13'b0000000010000: n5350 = n5349;
      13'b0000000001000: n5350 = n5349;
      13'b0000000000100: n5350 = n5349;
      13'b0000000000010: n5350 = n4971;
      13'b0000000000001: n5350 = n5349;
      default: n5350 = n5349;
    endcase
  assign n5351 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5352 = n5351;
      13'b0100000000000: n5352 = n5351;
      13'b0010000000000: n5352 = n5351;
      13'b0001000000000: n5352 = n5351;
      13'b0000100000000: n5352 = n5351;
      13'b0000010000000: n5352 = n5351;
      13'b0000001000000: n5352 = n5351;
      13'b0000000100000: n5352 = n5351;
      13'b0000000010000: n5352 = n5351;
      13'b0000000001000: n5352 = n5351;
      13'b0000000000100: n5352 = 1'b1;
      13'b0000000000010: n5352 = 1'b1;
      13'b0000000000001: n5352 = n5351;
      default: n5352 = n5351;
    endcase
  assign n5353 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5354 = n5353;
      13'b0100000000000: n5354 = n5353;
      13'b0010000000000: n5354 = n5353;
      13'b0001000000000: n5354 = n5353;
      13'b0000100000000: n5354 = n5353;
      13'b0000010000000: n5354 = n5353;
      13'b0000001000000: n5354 = n5353;
      13'b0000000100000: n5354 = n5353;
      13'b0000000010000: n5354 = n5353;
      13'b0000000001000: n5354 = n5353;
      13'b0000000000100: n5354 = n5353;
      13'b0000000000010: n5354 = n4973;
      13'b0000000000001: n5354 = n5353;
      default: n5354 = n5353;
    endcase
  assign n5355 = n1788[58:57]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5356 = n5355;
      13'b0100000000000: n5356 = n5355;
      13'b0010000000000: n5356 = n5230;
      13'b0001000000000: n5356 = n5214;
      13'b0000100000000: n5356 = n5355;
      13'b0000010000000: n5356 = n5355;
      13'b0000001000000: n5356 = n5355;
      13'b0000000100000: n5356 = n5355;
      13'b0000000010000: n5356 = n5355;
      13'b0000000001000: n5356 = n5355;
      13'b0000000000100: n5356 = n5355;
      13'b0000000000010: n5356 = n5355;
      13'b0000000000001: n5356 = n5355;
      default: n5356 = n5355;
    endcase
  assign n5357 = n1788[60:59]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5358 = n5357;
      13'b0100000000000: n5358 = n5357;
      13'b0010000000000: n5358 = n5357;
      13'b0001000000000: n5358 = n5357;
      13'b0000100000000: n5358 = n5180;
      13'b0000010000000: n5358 = n5357;
      13'b0000001000000: n5358 = n5357;
      13'b0000000100000: n5358 = n5357;
      13'b0000000010000: n5358 = n5357;
      13'b0000000001000: n5358 = n5357;
      13'b0000000000100: n5358 = n5357;
      13'b0000000000010: n5358 = n5357;
      13'b0000000000001: n5358 = n5357;
      default: n5358 = n5357;
    endcase
  assign n5359 = n5297[0]; // extract
  assign n5360 = n1896[0]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5361 = n5359;
      13'b0100000000000: n5361 = n5360;
      13'b0010000000000: n5361 = n5360;
      13'b0001000000000: n5361 = n5360;
      13'b0000100000000: n5361 = n5360;
      13'b0000010000000: n5361 = n5360;
      13'b0000001000000: n5361 = n5360;
      13'b0000000100000: n5361 = n5360;
      13'b0000000010000: n5361 = n5360;
      13'b0000000001000: n5361 = n5059;
      13'b0000000000100: n5361 = n5360;
      13'b0000000000010: n5361 = n5360;
      13'b0000000000001: n5361 = n5360;
      default: n5361 = n5360;
    endcase
  assign n5362 = n5297[1]; // extract
  assign n5363 = n1896[1]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5364 = n5362;
      13'b0100000000000: n5364 = n5363;
      13'b0010000000000: n5364 = n5363;
      13'b0001000000000: n5364 = n5363;
      13'b0000100000000: n5364 = n5363;
      13'b0000010000000: n5364 = n5363;
      13'b0000001000000: n5364 = n5363;
      13'b0000000100000: n5364 = n5363;
      13'b0000000010000: n5364 = n5094;
      13'b0000000001000: n5364 = n5363;
      13'b0000000000100: n5364 = n5363;
      13'b0000000000010: n5364 = n5363;
      13'b0000000000001: n5364 = n5363;
      default: n5364 = n5363;
    endcase
  assign n5365 = n1788[74]; // extract
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5366 = n5365;
      13'b0100000000000: n5366 = n5365;
      13'b0010000000000: n5366 = n5365;
      13'b0001000000000: n5366 = n5365;
      13'b0000100000000: n5366 = n5365;
      13'b0000010000000: n5366 = n5365;
      13'b0000001000000: n5366 = n5365;
      13'b0000000100000: n5366 = n5137;
      13'b0000000010000: n5366 = n5365;
      13'b0000000001000: n5366 = n5365;
      13'b0000000000100: n5366 = n5365;
      13'b0000000000010: n5366 = n5365;
      13'b0000000000001: n5366 = n5365;
      default: n5366 = n5365;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5368 = 1'b0;
      13'b0100000000000: n5368 = 1'b0;
      13'b0010000000000: n5368 = 1'b0;
      13'b0001000000000: n5368 = 1'b0;
      13'b0000100000000: n5368 = 1'b0;
      13'b0000010000000: n5368 = 1'b0;
      13'b0000001000000: n5368 = 1'b0;
      13'b0000000100000: n5368 = 1'b0;
      13'b0000000010000: n5368 = 1'b0;
      13'b0000000001000: n5368 = 1'b0;
      13'b0000000000100: n5368 = 1'b1;
      13'b0000000000010: n5368 = 1'b0;
      13'b0000000000001: n5368 = 1'b0;
      default: n5368 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5370 = 1'b0;
      13'b0100000000000: n5370 = 1'b0;
      13'b0010000000000: n5370 = 1'b0;
      13'b0001000000000: n5370 = 1'b0;
      13'b0000100000000: n5370 = 1'b0;
      13'b0000010000000: n5370 = 1'b0;
      13'b0000001000000: n5370 = 1'b0;
      13'b0000000100000: n5370 = 1'b0;
      13'b0000000010000: n5370 = 1'b0;
      13'b0000000001000: n5370 = 1'b0;
      13'b0000000000100: n5370 = 1'b0;
      13'b0000000000010: n5370 = 1'b1;
      13'b0000000000001: n5370 = 1'b0;
      default: n5370 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5372 = n5299;
      13'b0100000000000: n5372 = 2'b00;
      13'b0010000000000: n5372 = 2'b00;
      13'b0001000000000: n5372 = 2'b00;
      13'b0000100000000: n5372 = 2'b00;
      13'b0000010000000: n5372 = 2'b00;
      13'b0000001000000: n5372 = 2'b00;
      13'b0000000100000: n5372 = 2'b00;
      13'b0000000010000: n5372 = 2'b00;
      13'b0000000001000: n5372 = 2'b00;
      13'b0000000000100: n5372 = 2'b00;
      13'b0000000000010: n5372 = 2'b00;
      13'b0000000000001: n5372 = 2'b00;
      default: n5372 = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5374 = 1'b0;
      13'b0100000000000: n5374 = 1'b0;
      13'b0010000000000: n5374 = 1'b0;
      13'b0001000000000: n5374 = 1'b0;
      13'b0000100000000: n5374 = 1'b0;
      13'b0000010000000: n5374 = 1'b0;
      13'b0000001000000: n5374 = 1'b0;
      13'b0000000100000: n5374 = 1'b0;
      13'b0000000010000: n5374 = n5096;
      13'b0000000001000: n5374 = 1'b0;
      13'b0000000000100: n5374 = 1'b1;
      13'b0000000000010: n5374 = 1'b1;
      13'b0000000000001: n5374 = 1'b0;
      default: n5374 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5306)
      13'b1000000000000: n5375 = n5300;
      13'b0100000000000: n5375 = n2057;
      13'b0010000000000: n5375 = n5232;
      13'b0001000000000: n5375 = n5216;
      13'b0000100000000: n5375 = n5182;
      13'b0000010000000: n5375 = n2057;
      13'b0000001000000: n5375 = n2057;
      13'b0000000100000: n5375 = n2057;
      13'b0000000010000: n5375 = n2057;
      13'b0000000001000: n5375 = n2057;
      13'b0000000000100: n5375 = n5019;
      13'b0000000000010: n5375 = n4975;
      13'b0000000000001: n5375 = n2057;
      default: n5375 = n2057;
    endcase
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5376 = n4825 ? n4882 : n5307;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5377 = n4825 ? n4884 : n5312;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5378 = n4825 ? n4885 : n5313;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5379 = n4825 ? n2025 : n5314;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5380 = n4825 ? n2028 : n5315;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5381 = n4825 ? n4852 : n5316;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5383 = n4825 ? n4888 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5385 = n4825 ? n4891 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5387 = n4825 ? 1'b0 : n5318;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5389 = n4825 ? 1'b0 : n5320;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5390 = n4825 ? n1785 : n5321;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5391 = n4825 ? n2031 : n5322;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5392 = n4825 ? n4894 : n5325;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5394 = n4825 ? 1'b0 : n5327;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5396 = n4825 ? 1'b0 : n5330;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5398 = n4825 ? 1'b0 : n5332;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5399 = n4825 ? n4897 : n5336;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5401 = n4825 ? 1'b0 : n5338;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5403 = n4825 ? n4900 : 1'b0;
  assign n5404 = {n5350, n5348};
  assign n5405 = {n5358, n5356};
  assign n5406 = {n5364, n5361};
  assign n5407 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5408 = n4825 ? n5407 : n5340;
  assign n5409 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5410 = n4825 ? n5409 : n5342;
  assign n5411 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5412 = n4825 ? n5411 : n5344;
  assign n5413 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5414 = n4825 ? n5413 : n5346;
  assign n5415 = n5404[0]; // extract
  assign n5416 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5417 = n4825 ? n5416 : n5415;
  assign n5418 = n5404[1]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5419 = n4825 ? n4854 : n5418;
  assign n5420 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5421 = n4825 ? n5420 : n5352;
  assign n5422 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5423 = n4825 ? n5422 : n5354;
  assign n5424 = n1788[60:57]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5425 = n4825 ? n5424 : n5405;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5426 = n4838 & n4825;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5427 = n4825 ? n1896 : n5406;
  assign n5428 = n1788[74]; // extract
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5429 = n4825 ? n5428 : n5366;
  assign n5430 = {n5374, n5372};
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5432 = n4825 ? 1'b0 : n5368;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5434 = n4825 ? 1'b0 : n5370;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5436 = n4825 ? 3'b000 : n5430;
  /* TG68KdotC_Kernel.vhd:2420:57  */
  assign n5437 = n4825 ? n4905 : n5375;
  /* TG68KdotC_Kernel.vhd:2402:49  */
  assign n5439 = n3478 == 3'b111;
  assign n5440 = {n5439, n4824, n4714, n3943, n3803, n3696, n3597};
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5441 = n5376;
      7'b0100000: n5441 = make_berr;
      7'b0010000: n5441 = make_berr;
      7'b0001000: n5441 = make_berr;
      7'b0000100: n5441 = make_berr;
      7'b0000010: n5441 = n3677;
      7'b0000001: n5441 = n3508;
      default: n5441 = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5442 = n5377;
      7'b0100000: n5442 = n4804;
      7'b0010000: n5442 = n4636;
      7'b0001000: n5442 = n3848;
      7'b0000100: n5442 = n3725;
      7'b0000010: n5442 = n3625;
      7'b0000001: n5442 = n3517;
      default: n5442 = n1800;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5443 = n5378;
      7'b0100000: n5443 = n1903;
      7'b0010000: n5443 = n4637;
      7'b0001000: n5443 = n3846;
      7'b0000100: n5443 = n1903;
      7'b0000010: n5443 = n1903;
      7'b0000001: n5443 = n1903;
      default: n5443 = n1903;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5444 = n5379;
      7'b0100000: n5444 = n2025;
      7'b0010000: n5444 = n2025;
      7'b0001000: n5444 = n2025;
      7'b0000100: n5444 = n2025;
      7'b0000010: n5444 = n2025;
      7'b0000001: n5444 = n2025;
      default: n5444 = n2025;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5445 = n5380;
      7'b0100000: n5445 = n2028;
      7'b0010000: n5445 = n2028;
      7'b0001000: n5445 = n2028;
      7'b0000100: n5445 = n2028;
      7'b0000010: n5445 = n2028;
      7'b0000001: n5445 = n2028;
      default: n5445 = n2028;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5447 = 1'b0;
      7'b0100000: n5447 = n4806;
      7'b0010000: n5447 = n4639;
      7'b0001000: n5447 = n3924;
      7'b0000100: n5447 = n3787;
      7'b0000010: n5447 = n3680;
      7'b0000001: n5447 = n3573;
      default: n5447 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5448 = n5381;
      7'b0100000: n5448 = n1892;
      7'b0010000: n5448 = n4640;
      7'b0001000: n5448 = n1892;
      7'b0000100: n5448 = n1892;
      7'b0000010: n5448 = n1892;
      7'b0000001: n5448 = n1892;
      default: n5448 = n1892;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5450 = n5383;
      7'b0100000: n5450 = 1'b0;
      7'b0010000: n5450 = 1'b0;
      7'b0001000: n5450 = 1'b0;
      7'b0000100: n5450 = 1'b0;
      7'b0000010: n5450 = 1'b0;
      7'b0000001: n5450 = 1'b0;
      default: n5450 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5452 = 1'b0;
      7'b0100000: n5452 = n4808;
      7'b0010000: n5452 = 1'b0;
      7'b0001000: n5452 = 1'b0;
      7'b0000100: n5452 = 1'b0;
      7'b0000010: n5452 = 1'b0;
      7'b0000001: n5452 = 1'b0;
      default: n5452 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5454 = n5385;
      7'b0100000: n5454 = 1'b0;
      7'b0010000: n5454 = n4641;
      7'b0001000: n5454 = 1'b0;
      7'b0000100: n5454 = 1'b0;
      7'b0000010: n5454 = 1'b0;
      7'b0000001: n5454 = 1'b0;
      default: n5454 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5456 = n5387;
      7'b0100000: n5456 = n4810;
      7'b0010000: n5456 = n4643;
      7'b0001000: n5456 = 1'b0;
      7'b0000100: n5456 = 1'b0;
      7'b0000010: n5456 = 1'b0;
      7'b0000001: n5456 = 1'b0;
      default: n5456 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5458 = n5389;
      7'b0100000: n5458 = n4812;
      7'b0010000: n5458 = n4644;
      7'b0001000: n5458 = n3926;
      7'b0000100: n5458 = n3788;
      7'b0000010: n5458 = 1'b0;
      7'b0000001: n5458 = n3575;
      default: n5458 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5460 = 1'b0;
      7'b0100000: n5460 = 1'b0;
      7'b0010000: n5460 = n4646;
      7'b0001000: n5460 = 1'b0;
      7'b0000100: n5460 = 1'b0;
      7'b0000010: n5460 = 1'b0;
      7'b0000001: n5460 = 1'b0;
      default: n5460 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5462 = 1'b0;
      7'b0100000: n5462 = 1'b0;
      7'b0010000: n5462 = n4648;
      7'b0001000: n5462 = 1'b0;
      7'b0000100: n5462 = 1'b0;
      7'b0000010: n5462 = 1'b0;
      7'b0000001: n5462 = 1'b0;
      default: n5462 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5464 = 1'b0;
      7'b0100000: n5464 = 1'b0;
      7'b0010000: n5464 = n4650;
      7'b0001000: n5464 = 1'b0;
      7'b0000100: n5464 = 1'b0;
      7'b0000010: n5464 = 1'b0;
      7'b0000001: n5464 = 1'b0;
      default: n5464 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5465 = n5390;
      7'b0100000: n5465 = n1785;
      7'b0010000: n5465 = n1785;
      7'b0001000: n5465 = n1785;
      7'b0000100: n5465 = n1785;
      7'b0000010: n5465 = n1785;
      7'b0000001: n5465 = n1785;
      default: n5465 = n1785;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5467 = 1'b0;
      7'b0100000: n5467 = 1'b0;
      7'b0010000: n5467 = n4652;
      7'b0001000: n5467 = 1'b0;
      7'b0000100: n5467 = 1'b0;
      7'b0000010: n5467 = 1'b0;
      7'b0000001: n5467 = 1'b0;
      default: n5467 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5468 = n5391;
      7'b0100000: n5468 = n2031;
      7'b0010000: n5468 = n2031;
      7'b0001000: n5468 = n2031;
      7'b0000100: n5468 = n2031;
      7'b0000010: n5468 = n2031;
      7'b0000001: n5468 = n2031;
      default: n5468 = n2031;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5470 = n5392;
      7'b0100000: n5470 = n4814;
      7'b0010000: n5470 = n4653;
      7'b0001000: n5470 = n3927;
      7'b0000100: n5470 = n3789;
      7'b0000010: n5470 = n3682;
      7'b0000001: n5470 = n3578;
      default: n5470 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5472 = n5394;
      7'b0100000: n5472 = 1'b0;
      7'b0010000: n5472 = 1'b0;
      7'b0001000: n5472 = n3929;
      7'b0000100: n5472 = 1'b0;
      7'b0000010: n5472 = 1'b0;
      7'b0000001: n5472 = n3580;
      default: n5472 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5474 = n5396;
      7'b0100000: n5474 = 1'b0;
      7'b0010000: n5474 = 1'b0;
      7'b0001000: n5474 = 1'b0;
      7'b0000100: n5474 = 1'b0;
      7'b0000010: n5474 = 1'b0;
      7'b0000001: n5474 = 1'b0;
      default: n5474 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5476 = n5398;
      7'b0100000: n5476 = 1'b0;
      7'b0010000: n5476 = 1'b0;
      7'b0001000: n5476 = 1'b0;
      7'b0000100: n5476 = 1'b0;
      7'b0000010: n5476 = 1'b0;
      7'b0000001: n5476 = 1'b0;
      default: n5476 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5478 = n5399;
      7'b0100000: n5478 = n4816;
      7'b0010000: n5478 = n4654;
      7'b0001000: n5478 = n3930;
      7'b0000100: n5478 = n3790;
      7'b0000010: n5478 = n3684;
      7'b0000001: n5478 = n3582;
      default: n5478 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5480 = n5401;
      7'b0100000: n5480 = 1'b0;
      7'b0010000: n5480 = 1'b0;
      7'b0001000: n5480 = 1'b0;
      7'b0000100: n5480 = 1'b0;
      7'b0000010: n5480 = 1'b0;
      7'b0000001: n5480 = 1'b0;
      default: n5480 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5482 = n5403;
      7'b0100000: n5482 = n4818;
      7'b0010000: n5482 = n4656;
      7'b0001000: n5482 = n3931;
      7'b0000100: n5482 = n3791;
      7'b0000010: n5482 = n3686;
      7'b0000001: n5482 = n3584;
      default: n5482 = 1'b0;
    endcase
  assign n5483 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5484 = n5408;
      7'b0100000: n5484 = n5483;
      7'b0010000: n5484 = n4658;
      7'b0001000: n5484 = n5483;
      7'b0000100: n5484 = n5483;
      7'b0000010: n5484 = n5483;
      7'b0000001: n5484 = n5483;
      default: n5484 = n5483;
    endcase
  assign n5485 = n1788[20]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5486 = n5485;
      7'b0100000: n5486 = n5485;
      7'b0010000: n5486 = n4660;
      7'b0001000: n5486 = n5485;
      7'b0000100: n5486 = n5485;
      7'b0000010: n5486 = n5485;
      7'b0000001: n5486 = n5485;
      default: n5486 = n5485;
    endcase
  assign n5487 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5488 = n5410;
      7'b0100000: n5488 = n5487;
      7'b0010000: n5488 = n4662;
      7'b0001000: n5488 = n5487;
      7'b0000100: n5488 = n5487;
      7'b0000010: n5488 = n5487;
      7'b0000001: n5488 = n5487;
      default: n5488 = n5487;
    endcase
  assign n5489 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5490 = n5412;
      7'b0100000: n5490 = n5489;
      7'b0010000: n5490 = n4663;
      7'b0001000: n5490 = n5489;
      7'b0000100: n5490 = n5489;
      7'b0000010: n5490 = n5489;
      7'b0000001: n5490 = n5489;
      default: n5490 = n5489;
    endcase
  assign n5491 = n1788[36]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5492 = n5491;
      7'b0100000: n5492 = n5491;
      7'b0010000: n5492 = n4665;
      7'b0001000: n5492 = n5491;
      7'b0000100: n5492 = n5491;
      7'b0000010: n5492 = n5491;
      7'b0000001: n5492 = n5491;
      default: n5492 = n5491;
    endcase
  assign n5493 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5494 = n5493;
      7'b0100000: n5494 = n5493;
      7'b0010000: n5494 = n4667;
      7'b0001000: n5494 = n5493;
      7'b0000100: n5494 = n5493;
      7'b0000010: n5494 = n5493;
      7'b0000001: n5494 = n5493;
      default: n5494 = n5493;
    endcase
  assign n5495 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5496 = n5495;
      7'b0100000: n5496 = n5495;
      7'b0010000: n5496 = n4668;
      7'b0001000: n5496 = n5495;
      7'b0000100: n5496 = n5495;
      7'b0000010: n5496 = n5495;
      7'b0000001: n5496 = n5495;
      default: n5496 = n5495;
    endcase
  assign n5497 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5498 = n5414;
      7'b0100000: n5498 = n5497;
      7'b0010000: n5498 = n4670;
      7'b0001000: n5498 = n5497;
      7'b0000100: n5498 = n5497;
      7'b0000010: n5498 = n5497;
      7'b0000001: n5498 = n5497;
      default: n5498 = n5497;
    endcase
  assign n5499 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5500 = n5417;
      7'b0100000: n5500 = n5499;
      7'b0010000: n5500 = n5499;
      7'b0001000: n5500 = n5499;
      7'b0000100: n5500 = n5499;
      7'b0000010: n5500 = n5499;
      7'b0000001: n5500 = n5499;
      default: n5500 = n5499;
    endcase
  assign n5501 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5502 = n5419;
      7'b0100000: n5502 = n5501;
      7'b0010000: n5502 = n4672;
      7'b0001000: n5502 = n5501;
      7'b0000100: n5502 = n5501;
      7'b0000010: n5502 = n5501;
      7'b0000001: n5502 = n5501;
      default: n5502 = n5501;
    endcase
  assign n5503 = n1788[48]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5504 = n5503;
      7'b0100000: n5504 = n5503;
      7'b0010000: n5504 = n4675;
      7'b0001000: n5504 = n5503;
      7'b0000100: n5504 = n5503;
      7'b0000010: n5504 = n5503;
      7'b0000001: n5504 = n5503;
      default: n5504 = n5503;
    endcase
  assign n5505 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5506 = n5421;
      7'b0100000: n5506 = n5505;
      7'b0010000: n5506 = n4677;
      7'b0001000: n5506 = n5505;
      7'b0000100: n5506 = n5505;
      7'b0000010: n5506 = n5505;
      7'b0000001: n5506 = n5505;
      default: n5506 = n5505;
    endcase
  assign n5507 = n3832[0]; // extract
  assign n5508 = n1788[51]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5509 = n5508;
      7'b0100000: n5509 = n5508;
      7'b0010000: n5509 = n5508;
      7'b0001000: n5509 = n5507;
      7'b0000100: n5509 = n3723;
      7'b0000010: n5509 = n5508;
      7'b0000001: n5509 = n5508;
      default: n5509 = n5508;
    endcase
  assign n5510 = n3832[1]; // extract
  assign n5511 = n1788[52]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5512 = n5511;
      7'b0100000: n5512 = n5511;
      7'b0010000: n5512 = n5511;
      7'b0001000: n5512 = n5510;
      7'b0000100: n5512 = n5511;
      7'b0000010: n5512 = n5511;
      7'b0000001: n5512 = n5511;
      default: n5512 = n5511;
    endcase
  assign n5513 = n1788[53]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5514 = n5513;
      7'b0100000: n5514 = n5513;
      7'b0010000: n5514 = n5513;
      7'b0001000: n5514 = n3935;
      7'b0000100: n5514 = n5513;
      7'b0000010: n5514 = n5513;
      7'b0000001: n5514 = n5513;
      default: n5514 = n5513;
    endcase
  assign n5515 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5516 = n5515;
      7'b0100000: n5516 = n5515;
      7'b0010000: n5516 = n4680;
      7'b0001000: n5516 = n5515;
      7'b0000100: n5516 = n3795;
      7'b0000010: n5516 = n3688;
      7'b0000001: n5516 = n3586;
      default: n5516 = n5515;
    endcase
  assign n5517 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5518 = n5423;
      7'b0100000: n5518 = n5517;
      7'b0010000: n5518 = n4682;
      7'b0001000: n5518 = n5517;
      7'b0000100: n5518 = n5517;
      7'b0000010: n5518 = n5517;
      7'b0000001: n5518 = n5517;
      default: n5518 = n5517;
    endcase
  assign n5519 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5520 = n5519;
      7'b0100000: n5520 = n5519;
      7'b0010000: n5520 = n4685;
      7'b0001000: n5520 = n5519;
      7'b0000100: n5520 = n3797;
      7'b0000010: n5520 = n5519;
      7'b0000001: n5520 = n3588;
      default: n5520 = n5519;
    endcase
  assign n5521 = n1788[60:57]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5522 = n5425;
      7'b0100000: n5522 = n5521;
      7'b0010000: n5522 = n5521;
      7'b0001000: n5522 = n5521;
      7'b0000100: n5522 = n5521;
      7'b0000010: n5522 = n5521;
      7'b0000001: n5522 = n5521;
      default: n5522 = n5521;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5523 = n4904;
      7'b0100000: n5523 = n2055;
      7'b0010000: n5523 = n2055;
      7'b0001000: n5523 = n2055;
      7'b0000100: n5523 = n2055;
      7'b0000010: n5523 = n2055;
      7'b0000001: n5523 = n2055;
      default: n5523 = n2055;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5524 = n5427;
      7'b0100000: n5524 = n1896;
      7'b0010000: n5524 = n1896;
      7'b0001000: n5524 = n1896;
      7'b0000100: n5524 = n1896;
      7'b0000010: n5524 = n1896;
      7'b0000001: n5524 = n1896;
      default: n5524 = n1896;
    endcase
  assign n5525 = n1788[67]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5526 = n5525;
      7'b0100000: n5526 = n5525;
      7'b0010000: n5526 = n4687;
      7'b0001000: n5526 = n5525;
      7'b0000100: n5526 = n5525;
      7'b0000010: n5526 = n5525;
      7'b0000001: n5526 = n5525;
      default: n5526 = n5525;
    endcase
  assign n5527 = n1788[69]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5528 = n5527;
      7'b0100000: n5528 = n5527;
      7'b0010000: n5528 = n4689;
      7'b0001000: n5528 = n5527;
      7'b0000100: n5528 = n5527;
      7'b0000010: n5528 = n5527;
      7'b0000001: n5528 = n5527;
      default: n5528 = n5527;
    endcase
  assign n5529 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5530 = n5529;
      7'b0100000: n5530 = n5529;
      7'b0010000: n5530 = n4690;
      7'b0001000: n5530 = n5529;
      7'b0000100: n5530 = n5529;
      7'b0000010: n5530 = n5529;
      7'b0000001: n5530 = n5529;
      default: n5530 = n5529;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5531 = n2048;
      7'b0100000: n5531 = n2048;
      7'b0010000: n5531 = n4691;
      7'b0001000: n5531 = n2048;
      7'b0000100: n5531 = n2048;
      7'b0000010: n5531 = n2048;
      7'b0000001: n5531 = n2048;
      default: n5531 = n2048;
    endcase
  assign n5532 = n1788[74]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5533 = n5429;
      7'b0100000: n5533 = n5532;
      7'b0010000: n5533 = n5532;
      7'b0001000: n5533 = n5532;
      7'b0000100: n5533 = n5532;
      7'b0000010: n5533 = n5532;
      7'b0000001: n5533 = n5532;
      default: n5533 = n5532;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5535 = n5432;
      7'b0100000: n5535 = n4820;
      7'b0010000: n5535 = n4693;
      7'b0001000: n5535 = 1'b0;
      7'b0000100: n5535 = 1'b0;
      7'b0000010: n5535 = 1'b0;
      7'b0000001: n5535 = 1'b0;
      default: n5535 = 1'b0;
    endcase
  assign n5536 = n3591[0]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5538 = 1'b0;
      7'b0100000: n5538 = 1'b0;
      7'b0010000: n5538 = 1'b0;
      7'b0001000: n5538 = 1'b0;
      7'b0000100: n5538 = 1'b0;
      7'b0000010: n5538 = n3690;
      7'b0000001: n5538 = n5536;
      default: n5538 = 1'b0;
    endcase
  assign n5539 = n3591[1]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5541 = n5434;
      7'b0100000: n5541 = 1'b0;
      7'b0010000: n5541 = n4695;
      7'b0001000: n5541 = 1'b0;
      7'b0000100: n5541 = n3799;
      7'b0000010: n5541 = 1'b0;
      7'b0000001: n5541 = n5539;
      default: n5541 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5543 = 1'b0;
      7'b0100000: n5543 = 1'b0;
      7'b0010000: n5543 = 1'b0;
      7'b0001000: n5543 = 1'b0;
      7'b0000100: n5543 = 1'b0;
      7'b0000010: n5543 = n3692;
      7'b0000001: n5543 = 1'b0;
      default: n5543 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5545 = 1'b0;
      7'b0100000: n5545 = 1'b0;
      7'b0010000: n5545 = 1'b0;
      7'b0001000: n5545 = n3937;
      7'b0000100: n5545 = 1'b0;
      7'b0000010: n5545 = 1'b0;
      7'b0000001: n5545 = 1'b0;
      default: n5545 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5547 = 1'b0;
      7'b0100000: n5547 = 1'b0;
      7'b0010000: n5547 = n4697;
      7'b0001000: n5547 = 1'b0;
      7'b0000100: n5547 = 1'b0;
      7'b0000010: n5547 = 1'b0;
      7'b0000001: n5547 = 1'b0;
      default: n5547 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5549 = 1'b0;
      7'b0100000: n5549 = 1'b0;
      7'b0010000: n5549 = n4699;
      7'b0001000: n5549 = 1'b0;
      7'b0000100: n5549 = 1'b0;
      7'b0000010: n5549 = 1'b0;
      7'b0000001: n5549 = 1'b0;
      default: n5549 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5551 = 1'b0;
      7'b0100000: n5551 = 1'b0;
      7'b0010000: n5551 = n4701;
      7'b0001000: n5551 = 1'b0;
      7'b0000100: n5551 = 1'b0;
      7'b0000010: n5551 = 1'b0;
      7'b0000001: n5551 = 1'b0;
      default: n5551 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5553 = 1'b0;
      7'b0100000: n5553 = 1'b0;
      7'b0010000: n5553 = 1'b0;
      7'b0001000: n5553 = n3939;
      7'b0000100: n5553 = 1'b0;
      7'b0000010: n5553 = 1'b0;
      7'b0000001: n5553 = 1'b0;
      default: n5553 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5555 = 1'b0;
      7'b0100000: n5555 = 1'b0;
      7'b0010000: n5555 = n4703;
      7'b0001000: n5555 = 1'b0;
      7'b0000100: n5555 = 1'b0;
      7'b0000010: n5555 = 1'b0;
      7'b0000001: n5555 = n3593;
      default: n5555 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5557 = 1'b0;
      7'b0100000: n5557 = 1'b0;
      7'b0010000: n5557 = n4705;
      7'b0001000: n5557 = 1'b0;
      7'b0000100: n5557 = 1'b0;
      7'b0000010: n5557 = 1'b0;
      7'b0000001: n5557 = 1'b0;
      default: n5557 = 1'b0;
    endcase
  assign n5558 = n5436[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5560 = n5558;
      7'b0100000: n5560 = 2'b00;
      7'b0010000: n5560 = 2'b00;
      7'b0001000: n5560 = 2'b00;
      7'b0000100: n5560 = 2'b00;
      7'b0000010: n5560 = 2'b00;
      7'b0000001: n5560 = 2'b00;
      default: n5560 = 2'b00;
    endcase
  assign n5561 = n5436[2]; // extract
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5563 = n5561;
      7'b0100000: n5563 = n4822;
      7'b0010000: n5563 = n4706;
      7'b0001000: n5563 = n3941;
      7'b0000100: n5563 = n3801;
      7'b0000010: n5563 = n3694;
      7'b0000001: n5563 = n3595;
      default: n5563 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5565 = 1'b0;
      7'b0100000: n5565 = 1'b0;
      7'b0010000: n5565 = n4708;
      7'b0001000: n5565 = 1'b0;
      7'b0000100: n5565 = 1'b0;
      7'b0000010: n5565 = 1'b0;
      7'b0000001: n5565 = 1'b0;
      default: n5565 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5440)
      7'b1000000: n5566 = n5437;
      7'b0100000: n5566 = n2057;
      7'b0010000: n5566 = n4709;
      7'b0001000: n5566 = n2057;
      7'b0000100: n5566 = n2057;
      7'b0000010: n5566 = n2057;
      7'b0000001: n5566 = n2057;
      default: n5566 = n2057;
    endcase
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5567 = n3221 ? make_berr : n5441;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5568 = n3221 ? n3448 : n5442;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5569 = n3221 ? n3449 : n5443;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5570 = n3221 ? n2025 : n5444;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5571 = n3221 ? n2028 : n5445;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5573 = n3221 ? 1'b0 : n5447;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5574 = n3221 ? n1892 : n5448;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5576 = n3221 ? 1'b0 : n5450;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5578 = n3221 ? 1'b0 : n5452;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5579 = n3221 ? n3451 : n5454;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5580 = n3221 ? n3453 : n5456;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5581 = n3221 ? n3454 : n5458;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5583 = n3221 ? 1'b0 : n5460;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5585 = n3221 ? n3456 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5587 = n3221 ? 1'b0 : n5462;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5588 = n3221 ? n3457 : n5464;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5589 = n3221 ? n1785 : n5465;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5591 = n3221 ? 1'b0 : n5467;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5592 = n3221 ? n3458 : n5468;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5593 = n3221 ? n3459 : n5470;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5595 = n3221 ? 1'b0 : n5472;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5597 = n3221 ? 1'b0 : n5474;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5599 = n3221 ? 1'b0 : n5476;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5600 = n3221 ? n3460 : n5478;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5602 = n3221 ? 1'b0 : n5480;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5603 = n3221 ? n3461 : n5482;
  assign n5604 = {n5506, n5504, n5502, n5500};
  assign n5605 = {n5522, n5520, n5518, n5516, n5514, n5512, n5509};
  assign n5606 = {n5526, n5524, n5523};
  assign n5607 = {n5533, n5531};
  assign n5608 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5609 = n3221 ? n5608 : n5484;
  assign n5610 = n1788[20]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5611 = n3221 ? n5610 : n5486;
  assign n5612 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5613 = n3221 ? n5612 : n5488;
  assign n5614 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5615 = n3221 ? n5614 : n5490;
  assign n5616 = n1788[36]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5617 = n3221 ? n5616 : n5492;
  assign n5618 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5619 = n3221 ? n5618 : n5494;
  assign n5620 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5621 = n3221 ? n5620 : n5496;
  assign n5622 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5623 = n3221 ? n3463 : n5622;
  assign n5624 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5625 = n3221 ? n5624 : n5498;
  assign n5626 = n5604[2:0]; // extract
  assign n5627 = n1788[48]; // extract
  assign n5628 = {n5627, n2043};
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5629 = n3221 ? n5628 : n5626;
  assign n5630 = n5604[3]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5631 = n3221 ? n3465 : n5630;
  assign n5632 = n5605[4:0]; // extract
  assign n5633 = n1788[55:51]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5634 = n3221 ? n5633 : n5632;
  assign n5635 = n5605[5]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5636 = n3221 ? n3467 : n5635;
  assign n5637 = n5605[9:6]; // extract
  assign n5638 = n1788[60:57]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5639 = n3221 ? n5638 : n5637;
  assign n5640 = n1788[67]; // extract
  assign n5641 = {n5640, n1896, n2055};
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5642 = n3221 ? n5641 : n5606;
  assign n5643 = n1788[69]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5644 = n3221 ? n5643 : n5528;
  assign n5645 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5646 = n3221 ? n5645 : n5530;
  assign n5647 = n1788[74]; // extract
  assign n5648 = {n5647, n2048};
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5649 = n3221 ? n5648 : n5607;
  assign n5650 = {n5541, n5538};
  assign n5651 = {n5545, n5543};
  assign n5652 = {n5563, n5560};
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5653 = n3221 ? n3469 : n5535;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5655 = n3221 ? 2'b00 : n5650;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5657 = n3221 ? 2'b00 : n5651;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5658 = n3221 ? n3471 : n5547;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5660 = n3221 ? 1'b0 : n5549;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5662 = n3221 ? 1'b0 : n5551;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5664 = n3221 ? 1'b0 : n5553;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5666 = n3221 ? 1'b0 : n5555;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5668 = n3221 ? 1'b0 : n5557;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5670 = n3221 ? n3473 : 1'b0;
  assign n5671 = n5652[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5673 = n3221 ? 2'b00 : n5671;
  assign n5674 = n5652[2]; // extract
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5675 = n3221 ? n3475 : n5674;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5676 = n3221 ? n3477 : n5565;
  /* TG68KdotC_Kernel.vhd:1953:33  */
  assign n5677 = n3221 ? n2057 : n5566;
  /* TG68KdotC_Kernel.vhd:1952:25  */
  assign n5679 = n2058 == 4'b0100;
  /* TG68KdotC_Kernel.vhd:2631:50  */
  assign n5680 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2631:62  */
  assign n5682 = n5680 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2632:58  */
  assign n5683 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2632:70  */
  assign n5685 = n5683 == 3'b001;
  /* TG68KdotC_Kernel.vhd:2633:57  */
  assign n5689 = decodeopc ? 1'b1 : 1'b0;
  assign n5690 = n1788[53]; // extract
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5691 = n5886 ? 1'b1 : n5690;
  /* TG68KdotC_Kernel.vhd:2633:57  */
  assign n5693 = decodeopc ? 7'b0011001 : n2057;
  /* TG68KdotC_Kernel.vhd:2638:61  */
  assign n5694 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2638:73  */
  assign n5696 = n5694 == 3'b111;
  /* TG68KdotC_Kernel.vhd:2638:91  */
  assign n5697 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2638:103  */
  assign n5699 = n5697 == 2'b01;
  /* TG68KdotC_Kernel.vhd:2638:118  */
  assign n5700 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:2638:130  */
  assign n5702 = n5700 == 3'b100;
  /* TG68KdotC_Kernel.vhd:2638:109  */
  assign n5703 = n5699 | n5702;
  /* TG68KdotC_Kernel.vhd:2638:80  */
  assign n5704 = n5703 & n5696;
  /* TG68KdotC_Kernel.vhd:2639:63  */
  assign n5705 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:2640:74  */
  assign n5706 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2640:86  */
  assign n5708 = n5706 == 2'b01;
  /* TG68KdotC_Kernel.vhd:2642:90  */
  assign n5709 = opcode[0]; // extract
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5711 = n5790 ? 1'b1 : n2048;
  /* TG68KdotC_Kernel.vhd:2641:73  */
  assign n5712 = n5709 & decodeopc;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5714 = n5795 ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:2648:73  */
  assign n5716 = decodeopc ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2640:65  */
  assign n5717 = n5708 ? n1903 : n5716;
  /* TG68KdotC_Kernel.vhd:2640:65  */
  assign n5718 = n5712 & n5708;
  /* TG68KdotC_Kernel.vhd:2640:65  */
  assign n5719 = decodeopc & n5708;
  /* TG68KdotC_Kernel.vhd:2652:99  */
  assign n5720 = ~decodeopc;
  /* TG68KdotC_Kernel.vhd:2652:86  */
  assign n5721 = n5720 & exe_condition;
  /* TG68KdotC_Kernel.vhd:2652:65  */
  assign n5724 = n5721 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2652:65  */
  assign n5727 = n5721 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5728 = n5781 ? n5717 : n1903;
  /* TG68KdotC_Kernel.vhd:2639:57  */
  assign n5731 = n5705 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2639:57  */
  assign n5733 = n5705 ? n5724 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2639:57  */
  assign n5735 = n5705 ? n5727 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2639:57  */
  assign n5736 = n5718 & n5705;
  /* TG68KdotC_Kernel.vhd:2639:57  */
  assign n5737 = n5719 & n5705;
  /* TG68KdotC_Kernel.vhd:2660:62  */
  assign n5738 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2660:74  */
  assign n5740 = n5738 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2660:91  */
  assign n5741 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2660:103  */
  assign n5743 = n5741 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2660:82  */
  assign n5744 = n5740 | n5743;
  /* TG68KdotC_Kernel.vhd:2665:63  */
  assign n5746 = CPU[0]; // extract
  /* TG68KdotC_Kernel.vhd:2665:80  */
  assign n5748 = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2665:71  */
  assign n5749 = n5748 & n5746;
  /* TG68KdotC_Kernel.vhd:2665:99  */
  assign n5750 = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2665:86  */
  assign n5751 = n5750 & n5749;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5753 = n5760 ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2668:66  */
  assign n5754 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2668:78  */
  assign n5756 = n5754 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2668:57  */
  assign n5759 = n5756 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5760 = n5751 & n5744;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5762 = n5744 ? 2'b00 : n1800;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5765 = n5744 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5768 = n5744 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5771 = n5744 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5774 = n5744 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5776 = n5744 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2660:49  */
  assign n5778 = n5744 ? n5759 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5779 = n5704 ? make_berr : n5753;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5780 = n5704 ? n1800 : n5762;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5781 = n5705 & n5704;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5783 = n5704 ? 1'b0 : n5765;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5784 = n5704 ? n5731 : n5768;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5786 = n5704 ? n5733 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5787 = n5704 ? n5735 : n5771;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5789 = n5704 ? 1'b0 : n5774;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5790 = n5736 & n5704;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5792 = n5704 ? 1'b0 : n5776;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5794 = n5704 ? 1'b0 : n5778;
  /* TG68KdotC_Kernel.vhd:2638:49  */
  assign n5795 = n5737 & n5704;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5796 = n5685 ? make_berr : n5779;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5797 = n5685 ? n1800 : n5780;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5798 = n5685 ? n1903 : n5728;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5800 = n5685 ? n5689 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5802 = n5685 ? 1'b0 : n5783;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5804 = n5685 ? 1'b0 : n5784;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5806 = n5685 ? 1'b0 : n5786;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5808 = n5685 ? 1'b0 : n5787;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5810 = n5685 ? 1'b0 : n5789;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5812 = decodeopc & n5685;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5813 = n5685 ? n2048 : n5711;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5815 = n5685 ? 1'b0 : n5792;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5817 = n5685 ? 1'b0 : n5794;
  /* TG68KdotC_Kernel.vhd:2632:49  */
  assign n5818 = n5685 ? n5693 : n5714;
  /* TG68KdotC_Kernel.vhd:2676:58  */
  assign n5819 = opcode[7:3]; // extract
  /* TG68KdotC_Kernel.vhd:2676:70  */
  assign n5821 = n5819 != 5'b00001;
  /* TG68KdotC_Kernel.vhd:2677:59  */
  assign n5822 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2677:71  */
  assign n5824 = n5822 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2677:88  */
  assign n5825 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2677:100  */
  assign n5827 = n5825 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2677:79  */
  assign n5828 = n5824 | n5827;
  /* TG68KdotC_Kernel.vhd:2676:80  */
  assign n5829 = n5828 & n5821;
  /* TG68KdotC_Kernel.vhd:2679:66  */
  assign n5830 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2679:78  */
  assign n5832 = n5830 == 3'b001;
  assign n5834 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5835 = n5862 ? 1'b1 : n5834;
  /* TG68KdotC_Kernel.vhd:2682:66  */
  assign n5836 = opcode[8]; // extract
  assign n5838 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5839 = n5864 ? 1'b1 : n5838;
  /* TG68KdotC_Kernel.vhd:2689:66  */
  assign n5843 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2689:78  */
  assign n5845 = n5843 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2689:57  */
  assign n5848 = n5845 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5851 = n5829 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5854 = n5829 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5857 = n5829 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5860 = n5829 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5862 = n5832 & n5829;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5864 = n5836 & n5829;
  assign n5865 = {1'b1, 1'b1};
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5867 = n5829 ? n5865 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5869 = n5829 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2676:49  */
  assign n5871 = n5829 ? n5848 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5872 = n5682 ? n5796 : make_berr;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5873 = n5682 ? n5797 : n1800;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5874 = n5682 ? n5798 : n1903;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5876 = n5682 ? n5800 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5877 = n5682 ? n5802 : n5851;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5878 = n5682 ? n5804 : n5854;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5880 = n5682 ? n5806 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5881 = n5682 ? n5808 : n5857;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5882 = n5682 ? n5810 : n5860;
  assign n5883 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5884 = n5682 ? n5883 : n5835;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5886 = n5812 & n5682;
  assign n5887 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5888 = n5682 ? n5887 : n5839;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5889 = n5682 ? n5813 : n2048;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5891 = n5682 ? 2'b00 : n5867;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5893 = n5682 ? n5815 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5895 = n5682 ? 1'b0 : n5869;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5896 = n5682 ? n5817 : n5871;
  /* TG68KdotC_Kernel.vhd:2631:41  */
  assign n5897 = n5682 ? n5818 : n2057;
  /* TG68KdotC_Kernel.vhd:2630:25  */
  assign n5899 = n2058 == 4'b0101;
  /* TG68KdotC_Kernel.vhd:2702:47  */
  assign n5901 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2703:50  */
  assign n5902 = opcode[11:8]; // extract
  /* TG68KdotC_Kernel.vhd:2703:63  */
  assign n5904 = n5902 == 4'b0001;
  /* TG68KdotC_Kernel.vhd:2706:58  */
  assign n5906 = opcode[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:2706:70  */
  assign n5908 = n5906 == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:2709:61  */
  assign n5910 = opcode[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:2709:73  */
  assign n5912 = n5910 == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:2709:49  */
  assign n5914 = n5912 ? n1903 : 2'b11;
  /* TG68KdotC_Kernel.vhd:2709:49  */
  assign n5917 = n5912 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2709:49  */
  assign n5920 = n5912 ? 7'b0010111 : 7'b0010110;
  /* TG68KdotC_Kernel.vhd:2706:49  */
  assign n5921 = n5908 ? n1903 : n5914;
  /* TG68KdotC_Kernel.vhd:2706:49  */
  assign n5923 = n5908 ? 1'b0 : n5917;
  /* TG68KdotC_Kernel.vhd:2706:49  */
  assign n5924 = n5908 ? 1'b1 : n2048;
  /* TG68KdotC_Kernel.vhd:2706:49  */
  assign n5926 = n5908 ? 7'b0010111 : n5920;
  /* TG68KdotC_Kernel.vhd:2717:58  */
  assign n5927 = opcode[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:2717:70  */
  assign n5929 = n5927 == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:2720:61  */
  assign n5931 = opcode[7:0]; // extract
  /* TG68KdotC_Kernel.vhd:2720:73  */
  assign n5933 = n5931 == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:2720:49  */
  assign n5935 = n5933 ? n1903 : 2'b01;
  /* TG68KdotC_Kernel.vhd:2717:49  */
  assign n5936 = n5929 ? n1903 : n5935;
  /* TG68KdotC_Kernel.vhd:2717:49  */
  assign n5937 = n5929 ? 1'b1 : n2048;
  /* TG68KdotC_Kernel.vhd:2703:41  */
  assign n5938 = n5904 ? n5921 : n5936;
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5940 = n5949 ? 1'b1 : n1892;
  /* TG68KdotC_Kernel.vhd:2703:41  */
  assign n5942 = n5904 ? n5923 : 1'b0;
  assign n5943 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5944 = n5953 ? 1'b1 : n5943;
  /* TG68KdotC_Kernel.vhd:2703:41  */
  assign n5945 = n5904 ? n5924 : n5937;
  /* TG68KdotC_Kernel.vhd:2703:41  */
  assign n5947 = n5904 ? n5926 : 7'b0010101;
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5948 = n5901 ? n5938 : n1903;
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5949 = n5904 & n5901;
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5951 = n5901 ? n5942 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5953 = n5904 & n5901;
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5954 = n5901 ? n5945 : n2048;
  /* TG68KdotC_Kernel.vhd:2702:33  */
  assign n5955 = n5901 ? n5947 : n2057;
  /* TG68KdotC_Kernel.vhd:2699:25  */
  assign n5957 = n2058 == 4'b0110;
  /* TG68KdotC_Kernel.vhd:2731:42  */
  assign n5958 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2731:45  */
  assign n5959 = ~n5958;
  /* TG68KdotC_Kernel.vhd:2731:33  */
  assign n5964 = n5959 ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2731:33  */
  assign n5967 = n5959 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2731:33  */
  assign n5970 = n5959 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2731:33  */
  assign n5973 = n5959 ? 1'b0 : 1'b1;
  assign n5974 = {1'b1, 1'b1};
  /* TG68KdotC_Kernel.vhd:2731:33  */
  assign n5976 = n5959 ? n5974 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2731:33  */
  assign n5978 = n5959 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2730:25  */
  assign n5980 = n2058 == 4'b0111;
  /* TG68KdotC_Kernel.vhd:2744:42  */
  assign n5981 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2744:54  */
  assign n5983 = n5981 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2746:50  */
  assign n5984 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2746:62  */
  assign n5986 = n5984 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2745:56  */
  assign n5988 = n5986 & 1'b1;
  /* TG68KdotC_Kernel.vhd:2746:81  */
  assign n5989 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2746:93  */
  assign n5991 = n5989 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2746:111  */
  assign n5992 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2746:123  */
  assign n5994 = n5992 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2746:102  */
  assign n5995 = n5991 | n5994;
  /* TG68KdotC_Kernel.vhd:2746:70  */
  assign n5996 = n5995 & n5988;
  /* TG68KdotC_Kernel.vhd:2747:58  */
  assign n5997 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2747:70  */
  assign n5999 = n5997 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2747:49  */
  assign n6002 = n5999 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2750:64  */
  assign n6004 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2750:70  */
  assign n6005 = nextpass & n6004;
  /* TG68KdotC_Kernel.vhd:2750:98  */
  assign n6006 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2750:110  */
  assign n6008 = n6006 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2750:116  */
  assign n6009 = decodeopc & n6008;
  /* TG68KdotC_Kernel.vhd:2750:88  */
  assign n6010 = n6005 | n6009;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6012 = n6266 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6014 = n6050 ? 7'b1010101 : n2057;
  /* TG68KdotC_Kernel.vhd:2755:59  */
  assign n6015 = ~z_error;
  /* TG68KdotC_Kernel.vhd:2755:78  */
  assign n6016 = ~set_v_flag;
  /* TG68KdotC_Kernel.vhd:2755:64  */
  assign n6017 = n6016 & n6015;
  /* TG68KdotC_Kernel.vhd:2755:49  */
  assign n6020 = n6017 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2759:75  */
  assign n6021 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2759:87  */
  assign n6023 = n6021 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2759:93  */
  assign n6024 = decodeopc & n6023;
  /* TG68KdotC_Kernel.vhd:2759:65  */
  assign n6025 = nextpass | n6024;
  /* TG68KdotC_Kernel.vhd:2759:49  */
  assign n6028 = n6025 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6030 = n5996 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6031 = n6010 & n5996;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6033 = n5996 ? n6002 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6036 = n5996 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6038 = n5996 ? n6028 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6041 = n5996 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6044 = n5996 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6047 = n5996 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6049 = n5996 ? n6020 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2745:41  */
  assign n6050 = n6010 & n5996;
  /* TG68KdotC_Kernel.vhd:2767:45  */
  assign n6051 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2767:63  */
  assign n6052 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2767:75  */
  assign n6054 = n6052 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2767:53  */
  assign n6055 = n6054 & n6051;
  /* TG68KdotC_Kernel.vhd:2768:50  */
  assign n6056 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2768:62  */
  assign n6058 = n6056 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2773:53  */
  assign n6062 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2773:65  */
  assign n6064 = n6062 == 2'b01;
  /* TG68KdotC_Kernel.vhd:2773:80  */
  assign n6065 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2773:92  */
  assign n6067 = n6065 == 2'b10;
  /* TG68KdotC_Kernel.vhd:2773:71  */
  assign n6068 = n6064 | n6067;
  /* TG68KdotC_Kernel.vhd:2777:58  */
  assign n6071 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2777:71  */
  assign n6073 = n6071 == 2'b01;
  /* TG68KdotC_Kernel.vhd:2777:49  */
  assign n6078 = n6073 ? 2'b01 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2777:49  */
  assign n6080 = n6073 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2777:49  */
  assign n6082 = n6073 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2784:58  */
  assign n6083 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:2784:61  */
  assign n6084 = ~n6083;
  /* TG68KdotC_Kernel.vhd:2785:66  */
  assign n6085 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2785:79  */
  assign n6087 = n6085 == 2'b01;
  /* TG68KdotC_Kernel.vhd:2785:57  */
  assign n6090 = n6087 ? 2'b00 : 2'b01;
  assign n6094 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6095 = n6136 ? 1'b1 : n6094;
  assign n6096 = n1788[80]; // extract
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6097 = n6140 ? 1'b1 : n6096;
  /* TG68KdotC_Kernel.vhd:2792:57  */
  assign n6099 = decodeopc ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:2800:57  */
  assign n6101 = decodeopc ? 1'b1 : n2031;
  /* TG68KdotC_Kernel.vhd:2800:57  */
  assign n6103 = decodeopc ? 7'b0011110 : n2057;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6104 = n6120 ? n6090 : datatype;
  /* TG68KdotC_Kernel.vhd:2784:49  */
  assign n6107 = n6084 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2784:49  */
  assign n6110 = n6084 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2784:49  */
  assign n6111 = n6084 ? n2031 : n6101;
  /* TG68KdotC_Kernel.vhd:2784:49  */
  assign n6113 = decodeopc & n6084;
  /* TG68KdotC_Kernel.vhd:2784:49  */
  assign n6115 = decodeopc & n6084;
  /* TG68KdotC_Kernel.vhd:2784:49  */
  assign n6117 = n6084 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2784:49  */
  assign n6118 = n6084 ? n6099 : n6103;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6119 = n6068 ? n6078 : n1800;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6120 = n6084 & n6068;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6122 = n6068 ? n6107 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6125 = n6068 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6127 = n6068 ? n6110 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6128 = n6068 ? n6111 : n2031;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6131 = n6068 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6134 = n6068 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6136 = n6113 & n6068;
  assign n6137 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6138 = n6068 ? 1'b1 : n6137;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6140 = n6115 & n6068;
  assign n6141 = {n6082, n6080};
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6143 = n6068 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6145 = n6068 ? n6117 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6147 = n6068 ? n6141 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2773:41  */
  assign n6148 = n6068 ? n6118 : n2057;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6149 = n6058 ? n1800 : n6119;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6150 = n6058 ? datatype : n6104;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6152 = n6058 ? 1'b0 : n6122;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6154 = n6058 ? 1'b0 : n6125;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6156 = n6058 ? 1'b0 : n6127;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6157 = n6058 ? n2031 : n6128;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6159 = n6058 ? 1'b0 : n6131;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6161 = n6058 ? 1'b0 : n6134;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6164 = n6058 ? 1'b1 : 1'b0;
  assign n6165 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6166 = n6058 ? n6165 : n6095;
  assign n6167 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6168 = n6058 ? n6167 : n6138;
  assign n6169 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6170 = n6248 ? 1'b1 : n6169;
  assign n6171 = n1788[80]; // extract
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6172 = n6058 ? n6171 : n6097;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6174 = n6058 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6176 = n6058 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6178 = n6058 ? 1'b0 : n6143;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6180 = n6058 ? 1'b0 : n6145;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6182 = n6058 ? 2'b00 : n6147;
  /* TG68KdotC_Kernel.vhd:2768:41  */
  assign n6183 = n6058 ? n2057 : n6148;
  /* TG68KdotC_Kernel.vhd:2810:50  */
  assign n6184 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2810:62  */
  assign n6186 = n6184 != 2'b11;
  /* TG68KdotC_Kernel.vhd:2811:52  */
  assign n6187 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2811:55  */
  assign n6188 = ~n6187;
  /* TG68KdotC_Kernel.vhd:2811:70  */
  assign n6189 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2811:82  */
  assign n6191 = n6189 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2811:60  */
  assign n6192 = n6191 & n6188;
  /* TG68KdotC_Kernel.vhd:2811:101  */
  assign n6193 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2811:113  */
  assign n6195 = n6193 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2811:131  */
  assign n6196 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2811:143  */
  assign n6198 = n6196 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2811:122  */
  assign n6199 = n6195 | n6198;
  /* TG68KdotC_Kernel.vhd:2811:90  */
  assign n6200 = n6199 & n6192;
  /* TG68KdotC_Kernel.vhd:2812:51  */
  assign n6201 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2812:69  */
  assign n6202 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2812:81  */
  assign n6204 = n6202 != 2'b00;
  /* TG68KdotC_Kernel.vhd:2812:59  */
  assign n6205 = n6204 & n6201;
  /* TG68KdotC_Kernel.vhd:2812:99  */
  assign n6206 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2812:111  */
  assign n6208 = n6206 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2812:128  */
  assign n6209 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2812:140  */
  assign n6211 = n6209 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2812:119  */
  assign n6212 = n6208 | n6211;
  /* TG68KdotC_Kernel.vhd:2812:88  */
  assign n6213 = n6212 & n6205;
  /* TG68KdotC_Kernel.vhd:2811:151  */
  assign n6214 = n6200 | n6213;
  /* TG68KdotC_Kernel.vhd:2810:69  */
  assign n6215 = n6214 & n6186;
  /* TG68KdotC_Kernel.vhd:2810:41  */
  assign n6219 = n6215 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2810:41  */
  assign n6222 = n6215 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2810:41  */
  assign n6225 = n6215 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2810:41  */
  assign n6227 = n6215 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6228 = n6055 ? n6149 : n1800;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6229 = n6055 ? n6150 : datatype;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6231 = n6055 ? n6152 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6233 = n6055 ? n6154 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6235 = n6055 ? n6156 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6236 = n6055 ? n6157 : n2031;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6237 = n6055 ? n6159 : n6219;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6238 = n6055 ? n6161 : n6222;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6240 = n6055 ? 1'b0 : n6225;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6242 = n6055 ? n6164 : 1'b0;
  assign n6243 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6244 = n6055 ? n6166 : n6243;
  assign n6245 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6246 = n6055 ? n6168 : n6245;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6248 = n6058 & n6055;
  assign n6249 = n1788[80]; // extract
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6250 = n6055 ? n6172 : n6249;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6252 = n6055 ? n6174 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6254 = n6055 ? 1'b0 : n6227;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6256 = n6055 ? n6176 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6258 = n6055 ? n6178 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6260 = n6055 ? n6180 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6262 = n6055 ? n6182 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2767:33  */
  assign n6263 = n6055 ? n6183 : n2057;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6264 = n5983 ? n6030 : n6228;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6265 = n5983 ? datatype : n6229;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6266 = n6031 & n5983;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6268 = n5983 ? n6033 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6270 = n5983 ? 1'b0 : n6231;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6271 = n5983 ? n6036 : n6233;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6272 = n5983 ? n6038 : n6235;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6273 = n5983 ? n2031 : n6236;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6274 = n5983 ? n6041 : n6237;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6275 = n5983 ? n6044 : n6238;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6277 = n5983 ? n6047 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6279 = n5983 ? 1'b0 : n6240;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6281 = n5983 ? 1'b0 : n6242;
  assign n6282 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6283 = n5983 ? n6282 : n6244;
  assign n6284 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6285 = n5983 ? n6284 : n6246;
  assign n6286 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6287 = n5983 ? n6286 : n6170;
  assign n6288 = n1788[80]; // extract
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6289 = n5983 ? n6288 : n6250;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6291 = n5983 ? 1'b0 : n6252;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6293 = n5983 ? 1'b0 : n6254;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6295 = n5983 ? 1'b0 : n6256;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6297 = n5983 ? 1'b0 : n6258;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6298 = n5983 ? n6049 : n6260;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6300 = n5983 ? 2'b00 : n6262;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6301 = n5983 ? n6014 : n6263;
  /* TG68KdotC_Kernel.vhd:2743:25  */
  assign n6303 = n2058 == 4'b1000;
  /* TG68KdotC_Kernel.vhd:2823:42  */
  assign n6304 = opcode[8:3]; // extract
  /* TG68KdotC_Kernel.vhd:2823:54  */
  assign n6306 = n6304 != 6'b000001;
  /* TG68KdotC_Kernel.vhd:2824:45  */
  assign n6307 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2824:48  */
  assign n6308 = ~n6307;
  /* TG68KdotC_Kernel.vhd:2824:62  */
  assign n6309 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2824:74  */
  assign n6311 = n6309 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2824:53  */
  assign n6312 = n6308 | n6311;
  /* TG68KdotC_Kernel.vhd:2824:92  */
  assign n6313 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2824:104  */
  assign n6315 = n6313 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2824:122  */
  assign n6316 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2824:134  */
  assign n6318 = n6316 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2824:113  */
  assign n6319 = n6315 | n6318;
  /* TG68KdotC_Kernel.vhd:2824:81  */
  assign n6320 = n6319 & n6312;
  /* TG68KdotC_Kernel.vhd:2825:43  */
  assign n6321 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2825:62  */
  assign n6322 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2825:74  */
  assign n6324 = n6322 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2825:91  */
  assign n6325 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2825:103  */
  assign n6327 = n6325 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2825:82  */
  assign n6328 = n6324 | n6327;
  /* TG68KdotC_Kernel.vhd:2825:51  */
  assign n6329 = n6328 & n6321;
  /* TG68KdotC_Kernel.vhd:2824:142  */
  assign n6330 = n6320 | n6329;
  /* TG68KdotC_Kernel.vhd:2823:65  */
  assign n6331 = n6330 & n6306;
  /* TG68KdotC_Kernel.vhd:2828:50  */
  assign n6333 = opcode[14]; // extract
  /* TG68KdotC_Kernel.vhd:2828:54  */
  assign n6334 = ~n6333;
  assign n6336 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6337 = n6411 ? 1'b1 : n6336;
  /* TG68KdotC_Kernel.vhd:2831:50  */
  assign n6338 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2831:62  */
  assign n6340 = n6338 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2832:58  */
  assign n6341 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2832:61  */
  assign n6342 = ~n6341;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6344 = n6386 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2837:58  */
  assign n6346 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:2837:49  */
  assign n6349 = n6346 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2841:49  */
  assign n6353 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2841:49  */
  assign n6356 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2846:58  */
  assign n6357 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2846:76  */
  assign n6358 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2846:88  */
  assign n6360 = n6358 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2846:66  */
  assign n6361 = n6360 & n6357;
  /* TG68KdotC_Kernel.vhd:2846:49  */
  assign n6364 = n6361 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2846:49  */
  assign n6367 = n6361 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6368 = n6342 & n6340;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6370 = n6340 ? n6349 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6373 = n6340 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6375 = n6340 ? n6353 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6377 = n6340 ? n6356 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6379 = n6340 ? 1'b0 : n6364;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6381 = n6340 ? 1'b0 : n6367;
  assign n6382 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6383 = n6409 ? 1'b1 : n6382;
  /* TG68KdotC_Kernel.vhd:2831:41  */
  assign n6385 = n6340 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6386 = n6368 & n6331;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6388 = n6331 ? n6370 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6390 = n6331 ? n6373 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6392 = n6331 ? n6375 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6394 = n6331 ? n6377 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6397 = n6331 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6400 = n6331 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6403 = n6331 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6405 = n6331 ? n6379 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6407 = n6331 ? n6381 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6409 = n6340 & n6331;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6411 = n6334 & n6331;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6413 = n6331 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:33  */
  assign n6415 = n6331 ? n6385 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2822:25  */
  assign n6417 = n2058 == 4'b1001;
  /* TG68KdotC_Kernel.vhd:2822:36  */
  assign n6419 = n2058 == 4'b1101;
  /* TG68KdotC_Kernel.vhd:2822:36  */
  assign n6420 = n6417 | n6419;
  /* TG68KdotC_Kernel.vhd:2858:25  */
  assign n6422 = n2058 == 4'b1010;
  /* TG68KdotC_Kernel.vhd:2863:42  */
  assign n6423 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2863:54  */
  assign n6425 = n6423 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2864:50  */
  assign n6426 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2864:62  */
  assign n6428 = n6426 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2864:80  */
  assign n6429 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2864:92  */
  assign n6431 = n6429 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2864:71  */
  assign n6432 = n6428 | n6431;
  /* TG68KdotC_Kernel.vhd:2866:58  */
  assign n6433 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2866:61  */
  assign n6434 = ~n6433;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6437 = n6595 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2866:49  */
  assign n6439 = n6434 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2873:66  */
  assign n6441 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:2873:57  */
  assign n6444 = n6441 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2871:49  */
  assign n6446 = setexecopc ? n6444 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2871:49  */
  assign n6449 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2871:49  */
  assign n6452 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2871:49  */
  assign n6455 = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6457 = n6434 & n6432;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6459 = n6432 ? n6446 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6461 = n6432 ? n6449 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6463 = n6432 ? n6452 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6465 = n6432 ? n6455 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6468 = n6432 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6471 = n6432 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6474 = n6432 ? 1'b1 : 1'b0;
  assign n6475 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6476 = n6432 ? 1'b1 : n6475;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6478 = n6432 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2864:41  */
  assign n6480 = n6432 ? n6439 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2885:50  */
  assign n6481 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2886:58  */
  assign n6482 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2886:70  */
  assign n6484 = n6482 == 3'b001;
  /* TG68KdotC_Kernel.vhd:2890:74  */
  assign n6486 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:2890:86  */
  assign n6488 = n6486 == 3'b111;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6490 = n6584 ? 1'b1 : n2045;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6494 = n6576 ? 2'b10 : n1903;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6495 = n6581 ? 1'b1 : n1884;
  assign n6496 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6497 = n6583 ? 1'b1 : n6496;
  /* TG68KdotC_Kernel.vhd:2889:57  */
  assign n6498 = n6488 & decodeopc;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6500 = n6594 ? 7'b0100010 : n2057;
  /* TG68KdotC_Kernel.vhd:2901:66  */
  assign n6503 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2901:78  */
  assign n6505 = n6503 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2901:95  */
  assign n6506 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2901:107  */
  assign n6508 = n6506 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2901:86  */
  assign n6509 = n6505 | n6508;
  /* TG68KdotC_Kernel.vhd:2901:57  */
  assign n6513 = n6509 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2901:57  */
  assign n6516 = n6509 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2901:57  */
  assign n6519 = n6509 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2901:57  */
  assign n6522 = n6509 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2901:57  */
  assign n6524 = n6509 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6525 = decodeopc & n6484;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6527 = n6484 ? 1'b0 : n6513;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6529 = n6484 ? 1'b0 : n6516;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6531 = n6484 ? 1'b1 : n6519;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6533 = n6484 ? 1'b0 : n6522;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6534 = decodeopc & n6484;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6536 = decodeopc & n6484;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6537 = n6498 & n6484;
  assign n6538 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6539 = n6484 ? 1'b1 : n6538;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6541 = n6484 ? 1'b0 : n6524;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6543 = n6484 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6545 = n6484 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2886:49  */
  assign n6546 = decodeopc & n6484;
  /* TG68KdotC_Kernel.vhd:2911:58  */
  assign n6547 = opcode[8:3]; // extract
  /* TG68KdotC_Kernel.vhd:2911:70  */
  assign n6549 = n6547 != 6'b000001;
  /* TG68KdotC_Kernel.vhd:2912:59  */
  assign n6550 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2912:71  */
  assign n6552 = n6550 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2912:89  */
  assign n6553 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2912:101  */
  assign n6555 = n6553 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2912:80  */
  assign n6556 = n6552 | n6555;
  /* TG68KdotC_Kernel.vhd:2911:81  */
  assign n6557 = n6556 & n6549;
  /* TG68KdotC_Kernel.vhd:2911:49  */
  assign n6562 = n6557 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2911:49  */
  assign n6565 = n6557 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2911:49  */
  assign n6568 = n6557 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2911:49  */
  assign n6571 = n6557 ? 1'b1 : 1'b0;
  assign n6572 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:2911:49  */
  assign n6573 = n6557 ? 1'b1 : n6572;
  /* TG68KdotC_Kernel.vhd:2911:49  */
  assign n6575 = n6557 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6576 = n6525 & n6481;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6577 = n6481 ? n6527 : n6562;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6578 = n6481 ? n6529 : n6565;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6579 = n6481 ? n6531 : n6568;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6580 = n6481 ? n6533 : n6571;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6581 = n6534 & n6481;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6583 = n6536 & n6481;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6584 = n6537 & n6481;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6585 = n6481 ? n6539 : n6573;
  assign n6586 = {n6543, n6541};
  assign n6587 = n6586[0]; // extract
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6589 = n6481 ? n6587 : 1'b0;
  assign n6590 = n6586[1]; // extract
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6591 = n6481 ? n6590 : n6575;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6593 = n6481 ? n6545 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2885:41  */
  assign n6594 = n6546 & n6481;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6595 = n6457 & n6425;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6596 = n6425 ? n1903 : n6494;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6598 = n6425 ? n6459 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6600 = n6425 ? n6461 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6602 = n6425 ? n6463 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6604 = n6425 ? n6465 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6605 = n6425 ? n6468 : n6577;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6606 = n6425 ? n6471 : n6578;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6607 = n6425 ? n6474 : n6579;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6609 = n6425 ? 1'b0 : n6580;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6610 = n6425 ? n1884 : n6495;
  assign n6611 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6612 = n6425 ? n6611 : n6497;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6613 = n6425 ? n2045 : n6490;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6614 = n6425 ? n6476 : n6585;
  assign n6615 = {n6591, n6589};
  assign n6616 = n6615[0]; // extract
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6618 = n6425 ? 1'b0 : n6616;
  assign n6619 = n6615[1]; // extract
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6620 = n6425 ? n6478 : n6619;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6622 = n6425 ? n6480 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6624 = n6425 ? 1'b0 : n6593;
  /* TG68KdotC_Kernel.vhd:2863:33  */
  assign n6625 = n6425 ? n2057 : n6500;
  /* TG68KdotC_Kernel.vhd:2862:25  */
  assign n6627 = n2058 == 4'b1011;
  /* TG68KdotC_Kernel.vhd:2926:42  */
  assign n6628 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2926:54  */
  assign n6630 = n6628 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2928:50  */
  assign n6631 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2928:62  */
  assign n6633 = n6631 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2927:56  */
  assign n6635 = n6633 & 1'b1;
  /* TG68KdotC_Kernel.vhd:2928:81  */
  assign n6636 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2928:93  */
  assign n6638 = n6636 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2928:111  */
  assign n6639 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2928:123  */
  assign n6641 = n6639 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2928:102  */
  assign n6642 = n6638 | n6641;
  /* TG68KdotC_Kernel.vhd:2928:70  */
  assign n6643 = n6642 & n6635;
  /* TG68KdotC_Kernel.vhd:2929:58  */
  assign n6644 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2929:70  */
  assign n6646 = n6644 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2929:49  */
  assign n6649 = n6646 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2932:64  */
  assign n6651 = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2932:70  */
  assign n6652 = nextpass & n6651;
  /* TG68KdotC_Kernel.vhd:2932:98  */
  assign n6653 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2932:110  */
  assign n6655 = n6653 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2932:116  */
  assign n6656 = decodeopc & n6655;
  /* TG68KdotC_Kernel.vhd:2932:88  */
  assign n6657 = n6652 | n6656;
  /* TG68KdotC_Kernel.vhd:2932:49  */
  assign n6661 = n6657 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2932:49  */
  assign n6663 = n6657 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2945:77  */
  assign n6665 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2945:89  */
  assign n6667 = n6665 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2945:95  */
  assign n6668 = decodeopc & n6667;
  /* TG68KdotC_Kernel.vhd:2945:67  */
  assign n6669 = nextpass | n6668;
  /* TG68KdotC_Kernel.vhd:2945:49  */
  assign n6672 = n6669 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2949:49  */
  assign n6675 = setexecopc ? 2'b10 : 2'b01;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6677 = n6643 ? n6675 : n1800;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6679 = n6643 ? n6649 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6682 = n6643 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6684 = n6643 ? n6672 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6687 = n6643 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6690 = n6643 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6693 = n6643 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6695 = n6643 ? n6661 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6697 = n6643 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2927:41  */
  assign n6699 = n6643 ? n6663 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2956:45  */
  assign n6700 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2956:63  */
  assign n6701 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2956:75  */
  assign n6703 = n6701 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2956:53  */
  assign n6704 = n6703 & n6700;
  /* TG68KdotC_Kernel.vhd:2957:50  */
  assign n6705 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2957:62  */
  assign n6707 = n6705 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2962:58  */
  assign n6710 = opcode[7:4]; // extract
  /* TG68KdotC_Kernel.vhd:2962:70  */
  assign n6712 = n6710 == 4'b0100;
  /* TG68KdotC_Kernel.vhd:2962:87  */
  assign n6713 = opcode[7:3]; // extract
  /* TG68KdotC_Kernel.vhd:2962:99  */
  assign n6715 = n6713 == 5'b10001;
  /* TG68KdotC_Kernel.vhd:2962:78  */
  assign n6716 = n6712 | n6715;
  /* TG68KdotC_Kernel.vhd:2967:66  */
  assign n6720 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:2967:84  */
  assign n6721 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:2967:74  */
  assign n6722 = n6721 & n6720;
  /* TG68KdotC_Kernel.vhd:2967:57  */
  assign n6725 = n6722 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2967:57  */
  assign n6728 = n6722 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6730 = n6736 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:2971:57  */
  assign n6733 = decodeopc ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6735 = n6716 ? 2'b10 : n1800;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6736 = decodeopc & n6716;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6738 = n6716 ? n6725 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6740 = n6716 ? n6728 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6742 = n6716 ? n6733 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6745 = n6716 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6748 = n6716 ? 1'b0 : 1'b1;
  assign n6749 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6750 = n6716 ? 1'b1 : n6749;
  assign n6751 = n1788[61]; // extract
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6752 = n6716 ? 1'b1 : n6751;
  assign n6753 = n1788[85]; // extract
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6754 = n6716 ? 1'b1 : n6753;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6755 = n6707 ? n1800 : n6735;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6756 = n6707 ? n1903 : n6730;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6758 = n6707 ? 1'b0 : n6738;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6760 = n6707 ? 1'b0 : n6740;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6762 = n6707 ? 1'b0 : n6742;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6764 = n6707 ? 1'b0 : n6745;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6766 = n6707 ? 1'b0 : n6748;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6769 = n6707 ? 1'b1 : 1'b0;
  assign n6770 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6771 = n6707 ? n6770 : n6750;
  assign n6772 = n1788[61]; // extract
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6773 = n6707 ? n6772 : n6752;
  assign n6774 = n1788[85]; // extract
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6775 = n6707 ? n6774 : n6754;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6777 = n6707 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2957:41  */
  assign n6779 = n6707 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2982:50  */
  assign n6780 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2982:62  */
  assign n6782 = n6780 != 2'b11;
  /* TG68KdotC_Kernel.vhd:2983:52  */
  assign n6783 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2983:55  */
  assign n6784 = ~n6783;
  /* TG68KdotC_Kernel.vhd:2983:70  */
  assign n6785 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2983:82  */
  assign n6787 = n6785 != 3'b001;
  /* TG68KdotC_Kernel.vhd:2983:60  */
  assign n6788 = n6787 & n6784;
  /* TG68KdotC_Kernel.vhd:2983:101  */
  assign n6789 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:2983:113  */
  assign n6791 = n6789 != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2983:131  */
  assign n6792 = opcode[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:2983:143  */
  assign n6794 = n6792 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2983:122  */
  assign n6795 = n6791 | n6794;
  /* TG68KdotC_Kernel.vhd:2983:90  */
  assign n6796 = n6795 & n6788;
  /* TG68KdotC_Kernel.vhd:2984:51  */
  assign n6797 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:2984:69  */
  assign n6798 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2984:81  */
  assign n6800 = n6798 != 2'b00;
  /* TG68KdotC_Kernel.vhd:2984:59  */
  assign n6801 = n6800 & n6797;
  /* TG68KdotC_Kernel.vhd:2984:99  */
  assign n6802 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2984:111  */
  assign n6804 = n6802 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2984:128  */
  assign n6805 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2984:140  */
  assign n6807 = n6805 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2984:119  */
  assign n6808 = n6804 | n6807;
  /* TG68KdotC_Kernel.vhd:2984:88  */
  assign n6809 = n6808 & n6801;
  /* TG68KdotC_Kernel.vhd:2983:151  */
  assign n6810 = n6796 | n6809;
  /* TG68KdotC_Kernel.vhd:2982:69  */
  assign n6811 = n6810 & n6782;
  /* TG68KdotC_Kernel.vhd:2982:41  */
  assign n6815 = n6811 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2982:41  */
  assign n6818 = n6811 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2982:41  */
  assign n6821 = n6811 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2982:41  */
  assign n6823 = n6811 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6824 = n6704 ? n6755 : n1800;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6825 = n6704 ? n6756 : n1903;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6827 = n6704 ? n6758 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6829 = n6704 ? n6760 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6831 = n6704 ? n6762 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6832 = n6704 ? n6764 : n6815;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6833 = n6704 ? n6766 : n6818;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6835 = n6704 ? 1'b0 : n6821;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6837 = n6704 ? n6769 : 1'b0;
  assign n6838 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6839 = n6704 ? n6771 : n6838;
  assign n6840 = n1788[61]; // extract
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6841 = n6704 ? n6773 : n6840;
  assign n6842 = n1788[85]; // extract
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6843 = n6704 ? n6775 : n6842;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6845 = n6704 ? n6777 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6847 = n6704 ? 1'b0 : n6823;
  /* TG68KdotC_Kernel.vhd:2956:33  */
  assign n6849 = n6704 ? n6779 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6850 = n6630 ? n6677 : n6824;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6851 = n6630 ? n1903 : n6825;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6853 = n6630 ? n6679 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6855 = n6630 ? 1'b0 : n6827;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6857 = n6630 ? n6682 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6859 = n6630 ? 1'b0 : n6829;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6860 = n6630 ? n6684 : n6831;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6861 = n6630 ? n6687 : n6832;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6862 = n6630 ? n6690 : n6833;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6864 = n6630 ? n6693 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6866 = n6630 ? 1'b0 : n6835;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6868 = n6630 ? 1'b0 : n6837;
  assign n6869 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6870 = n6630 ? n6869 : n6839;
  assign n6871 = n1788[61]; // extract
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6872 = n6630 ? n6871 : n6841;
  assign n6873 = n1788[85]; // extract
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6874 = n6630 ? n6873 : n6843;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6876 = n6630 ? 1'b0 : n6845;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6878 = n6630 ? 1'b0 : n6847;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6880 = n6630 ? 1'b0 : n6849;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6882 = n6630 ? n6695 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6884 = n6630 ? n6697 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2926:33  */
  assign n6886 = n6630 ? n6699 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2925:25  */
  assign n6888 = n2058 == 4'b1100;
  /* TG68KdotC_Kernel.vhd:2995:42  */
  assign n6889 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:2995:54  */
  assign n6891 = n6889 == 2'b11;
  /* TG68KdotC_Kernel.vhd:2996:50  */
  assign n6892 = opcode[11]; // extract
  /* TG68KdotC_Kernel.vhd:2996:54  */
  assign n6893 = ~n6892;
  /* TG68KdotC_Kernel.vhd:2997:54  */
  assign n6894 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:2997:66  */
  assign n6896 = n6894 != 2'b00;
  /* TG68KdotC_Kernel.vhd:2997:84  */
  assign n6897 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:2997:96  */
  assign n6899 = n6897 != 3'b111;
  /* TG68KdotC_Kernel.vhd:2997:113  */
  assign n6900 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:2997:125  */
  assign n6902 = n6900 == 2'b00;
  /* TG68KdotC_Kernel.vhd:2997:104  */
  assign n6903 = n6899 | n6902;
  /* TG68KdotC_Kernel.vhd:2997:73  */
  assign n6904 = n6903 & n6896;
  /* TG68KdotC_Kernel.vhd:3005:79  */
  assign n6906 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n6909 = n7237 ? 2'b01 : n1800;
  /* TG68KdotC_Kernel.vhd:2997:44  */
  assign n6912 = n6904 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n6913 = n7168 ? n6906 : n1779;
  /* TG68KdotC_Kernel.vhd:2997:44  */
  assign n6916 = n6904 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2997:44  */
  assign n6919 = n6904 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2997:44  */
  assign n6922 = n6904 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2997:44  */
  assign n6924 = n6904 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2997:44  */
  assign n6926 = n6904 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3013:70  */
  assign n6927 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3013:73  */
  assign n6928 = ~n6927;
  /* TG68KdotC_Kernel.vhd:3013:78  */
  assign n6930 = 1'b1 & n6928;
  /* TG68KdotC_Kernel.vhd:3013:63  */
  assign n6932 = 1'b0 | n6930;
  /* TG68KdotC_Kernel.vhd:3014:60  */
  assign n6933 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:3014:73  */
  assign n6935 = n6933 == 2'b11;
  /* TG68KdotC_Kernel.vhd:3014:88  */
  assign n6936 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3014:101  */
  assign n6938 = n6936 == 3'b010;
  /* TG68KdotC_Kernel.vhd:3014:79  */
  assign n6939 = n6935 | n6938;
  /* TG68KdotC_Kernel.vhd:3014:117  */
  assign n6940 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3014:130  */
  assign n6942 = n6940 == 3'b100;
  /* TG68KdotC_Kernel.vhd:3014:108  */
  assign n6943 = n6939 | n6942;
  /* TG68KdotC_Kernel.vhd:3015:59  */
  assign n6944 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3015:71  */
  assign n6946 = n6944 == 3'b001;
  /* TG68KdotC_Kernel.vhd:3015:87  */
  assign n6947 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3015:99  */
  assign n6949 = n6947 == 3'b011;
  /* TG68KdotC_Kernel.vhd:3015:78  */
  assign n6950 = n6946 | n6949;
  /* TG68KdotC_Kernel.vhd:3015:115  */
  assign n6951 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3015:127  */
  assign n6953 = n6951 == 3'b100;
  /* TG68KdotC_Kernel.vhd:3015:106  */
  assign n6954 = n6950 | n6953;
  /* TG68KdotC_Kernel.vhd:3015:144  */
  assign n6955 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3015:156  */
  assign n6957 = n6955 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3015:173  */
  assign n6958 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:3015:185  */
  assign n6960 = n6958 != 2'b00;
  /* TG68KdotC_Kernel.vhd:3015:163  */
  assign n6961 = n6960 & n6957;
  /* TG68KdotC_Kernel.vhd:3015:134  */
  assign n6962 = n6954 | n6961;
  /* TG68KdotC_Kernel.vhd:3014:138  */
  assign n6963 = n6962 & n6943;
  /* TG68KdotC_Kernel.vhd:3013:94  */
  assign n6964 = n6932 | n6963;
  /* TG68KdotC_Kernel.vhd:3016:60  */
  assign n6965 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:3016:73  */
  assign n6967 = n6965 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3016:88  */
  assign n6968 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3016:101  */
  assign n6970 = n6968 == 3'b011;
  /* TG68KdotC_Kernel.vhd:3016:79  */
  assign n6971 = n6967 | n6970;
  /* TG68KdotC_Kernel.vhd:3016:117  */
  assign n6972 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3016:130  */
  assign n6974 = n6972 == 3'b101;
  /* TG68KdotC_Kernel.vhd:3016:108  */
  assign n6975 = n6971 | n6974;
  /* TG68KdotC_Kernel.vhd:3017:59  */
  assign n6976 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3017:71  */
  assign n6978 = n6976 == 3'b001;
  /* TG68KdotC_Kernel.vhd:3017:87  */
  assign n6979 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3017:99  */
  assign n6981 = n6979 == 3'b011;
  /* TG68KdotC_Kernel.vhd:3017:78  */
  assign n6982 = n6978 | n6981;
  /* TG68KdotC_Kernel.vhd:3017:115  */
  assign n6983 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3017:127  */
  assign n6985 = n6983 == 3'b100;
  /* TG68KdotC_Kernel.vhd:3017:106  */
  assign n6986 = n6982 | n6985;
  /* TG68KdotC_Kernel.vhd:3017:143  */
  assign n6987 = opcode[5:2]; // extract
  /* TG68KdotC_Kernel.vhd:3017:155  */
  assign n6989 = n6987 == 4'b1111;
  /* TG68KdotC_Kernel.vhd:3017:134  */
  assign n6990 = n6986 | n6989;
  /* TG68KdotC_Kernel.vhd:3016:138  */
  assign n6991 = n6990 & n6975;
  /* TG68KdotC_Kernel.vhd:3015:195  */
  assign n6992 = n6964 | n6991;
  assign n6995 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:3021:57  */
  assign n6996 = decodeopc ? 1'b1 : n6995;
  assign n6997 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:3021:57  */
  assign n6998 = decodeopc ? 1'b1 : n6997;
  /* TG68KdotC_Kernel.vhd:3021:57  */
  assign n7000 = decodeopc ? 7'b0000001 : n2057;
  /* TG68KdotC_Kernel.vhd:3028:66  */
  assign n7002 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:3028:84  */
  assign n7003 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:3028:87  */
  assign n7004 = ~n7003;
  /* TG68KdotC_Kernel.vhd:3028:75  */
  assign n7005 = n7002 | n7004;
  /* TG68KdotC_Kernel.vhd:3028:57  */
  assign n7008 = n7005 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3031:66  */
  assign n7009 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3031:79  */
  assign n7011 = n7009 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3031:57  */
  assign n7014 = n7011 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3034:66  */
  assign n7015 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3034:79  */
  assign n7017 = n7015 == 3'b010;
  /* TG68KdotC_Kernel.vhd:3034:95  */
  assign n7018 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3034:108  */
  assign n7020 = n7018 == 3'b100;
  /* TG68KdotC_Kernel.vhd:3034:86  */
  assign n7021 = n7017 | n7020;
  /* TG68KdotC_Kernel.vhd:3034:124  */
  assign n7022 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3034:137  */
  assign n7024 = n7022 == 3'b110;
  /* TG68KdotC_Kernel.vhd:3034:115  */
  assign n7025 = n7021 | n7024;
  /* TG68KdotC_Kernel.vhd:3034:153  */
  assign n7026 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3034:166  */
  assign n7028 = n7026 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3034:144  */
  assign n7029 = n7025 | n7028;
  /* TG68KdotC_Kernel.vhd:3034:57  */
  assign n7032 = n7029 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3038:66  */
  assign n7033 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3038:79  */
  assign n7035 = n7033 == 3'b001;
  /* TG68KdotC_Kernel.vhd:3038:95  */
  assign n7036 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3038:108  */
  assign n7038 = n7036 == 3'b011;
  /* TG68KdotC_Kernel.vhd:3038:86  */
  assign n7039 = n7035 | n7038;
  /* TG68KdotC_Kernel.vhd:3038:124  */
  assign n7040 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3038:137  */
  assign n7042 = n7040 == 3'b101;
  /* TG68KdotC_Kernel.vhd:3038:115  */
  assign n7043 = n7039 | n7042;
  /* TG68KdotC_Kernel.vhd:3038:57  */
  assign n7046 = n7043 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3041:66  */
  assign n7047 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:3041:78  */
  assign n7049 = n7047 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3042:74  */
  assign n7050 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3042:87  */
  assign n7052 = n7050 != 3'b000;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7054 = n7074 ? 1'b1 : n7046;
  /* TG68KdotC_Kernel.vhd:3045:72  */
  assign n7055 = exec[42]; // extract
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7058 = n7067 ? 2'b01 : n1903;
  /* TG68KdotC_Kernel.vhd:3045:65  */
  assign n7061 = n7055 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3045:65  */
  assign n7064 = n7055 ? 1'b1 : 1'b0;
  assign n7065 = n1788[29]; // extract
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7066 = n7073 ? 1'b1 : n7065;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7067 = n7055 & n7049;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7069 = n7049 ? n7061 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7071 = n7049 ? n7064 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7073 = n7055 & n7049;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7074 = n7052 & n7049;
  /* TG68KdotC_Kernel.vhd:3052:63  */
  assign n7075 = set[62]; // extract
  /* TG68KdotC_Kernel.vhd:3052:57  */
  assign n7077 = n7075 ? 2'b01 : n7058;
  /* TG68KdotC_Kernel.vhd:3055:64  */
  assign n7078 = exec[62]; // extract
  /* TG68KdotC_Kernel.vhd:3055:57  */
  assign n7082 = n7078 ? 2'b01 : n7077;
  /* TG68KdotC_Kernel.vhd:3055:57  */
  assign n7084 = n7078 ? 1'b1 : n7069;
  /* TG68KdotC_Kernel.vhd:3055:57  */
  assign n7086 = n7078 ? 1'b1 : n7071;
  /* TG68KdotC_Kernel.vhd:3055:57  */
  assign n7087 = n7078 ? 1'b1 : n7066;
  assign n7088 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:3055:57  */
  assign n7089 = n7078 ? 1'b1 : n7088;
  /* TG68KdotC_Kernel.vhd:3055:57  */
  assign n7091 = n7078 ? 7'b1010000 : n7000;
  /* TG68KdotC_Kernel.vhd:3064:74  */
  assign n7092 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3064:87  */
  assign n7094 = n7092 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3064:65  */
  assign n7097 = n7094 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3064:65  */
  assign n7100 = n7094 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3069:74  */
  assign n7101 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3069:87  */
  assign n7103 = n7101 == 3'b001;
  /* TG68KdotC_Kernel.vhd:3069:103  */
  assign n7104 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3069:116  */
  assign n7106 = n7104 == 3'b011;
  /* TG68KdotC_Kernel.vhd:3069:94  */
  assign n7107 = n7103 | n7106;
  /* TG68KdotC_Kernel.vhd:3069:132  */
  assign n7108 = opcode[10:8]; // extract
  /* TG68KdotC_Kernel.vhd:3069:145  */
  assign n7110 = n7108 == 3'b101;
  /* TG68KdotC_Kernel.vhd:3069:123  */
  assign n7111 = n7107 | n7110;
  /* TG68KdotC_Kernel.vhd:3063:57  */
  assign n7113 = n7118 ? 1'b1 : n7086;
  /* TG68KdotC_Kernel.vhd:3063:57  */
  assign n7115 = setexecopc ? n7097 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3063:57  */
  assign n7117 = setexecopc ? n7100 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3063:57  */
  assign n7118 = n7111 & setexecopc;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7119 = n6992 ? n1903 : n7082;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7121 = n6992 ? 1'b0 : n7032;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7124 = n6992 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7126 = n6992 ? 1'b0 : n7115;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7128 = n6992 ? 1'b0 : n7117;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7130 = n6992 ? 1'b0 : n7084;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7132 = n6992 ? 1'b0 : n7113;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7135 = n6992 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7138 = n6992 ? 1'b1 : 1'b0;
  assign n7139 = n1788[29]; // extract
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7140 = n6992 ? n7139 : n7087;
  assign n7141 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7142 = n6992 ? n7141 : n6996;
  assign n7143 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7144 = n6992 ? n7143 : n7089;
  assign n7145 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7146 = n6992 ? n7145 : n6998;
  assign n7147 = {n7008, 1'b1};
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7149 = n6992 ? 1'b0 : n7014;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7151 = n6992 ? 1'b0 : n7054;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7153 = n6992 ? 2'b00 : n7147;
  /* TG68KdotC_Kernel.vhd:3013:49  */
  assign n7154 = n6992 ? n2057 : n7091;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7155 = n6904 & n6893;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7156 = n6893 ? n1903 : n7119;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7157 = n6893 ? n6912 : n7121;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7159 = n6893 ? 1'b0 : n7124;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7161 = n6893 ? 1'b0 : n7126;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7163 = n6893 ? 1'b0 : n7128;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7165 = n6893 ? 1'b0 : n7130;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7167 = n6893 ? 1'b0 : n7132;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7168 = n6904 & n6893;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7169 = n6893 ? n6916 : n7135;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7170 = n6893 ? n6919 : n7138;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7172 = n6893 ? n6922 : 1'b0;
  assign n7173 = n1788[29]; // extract
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7174 = n6893 ? n7173 : n7140;
  assign n7175 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7176 = n6893 ? n7175 : n7142;
  assign n7177 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7178 = n6893 ? n7177 : n7144;
  assign n7179 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7180 = n6893 ? n7179 : n7146;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7181 = n6893 ? n6924 : n7149;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7183 = n6893 ? 1'b0 : n7151;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7185 = n6893 ? 2'b00 : n7153;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7187 = n6893 ? n6926 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2996:41  */
  assign n7188 = n6893 ? n2057 : n7154;
  /* TG68KdotC_Kernel.vhd:3077:67  */
  assign n7189 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3077:70  */
  assign n7190 = ~n7189;
  /* TG68KdotC_Kernel.vhd:3077:75  */
  assign n7192 = 1'b1 & n7190;
  /* TG68KdotC_Kernel.vhd:3077:60  */
  assign n7194 = 1'b0 | n7192;
  /* TG68KdotC_Kernel.vhd:3079:71  */
  assign n7196 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:3082:66  */
  assign n7198 = opcode[5]; // extract
  /* TG68KdotC_Kernel.vhd:3087:98  */
  assign n7200 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3088:74  */
  assign n7201 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3088:87  */
  assign n7203 = n7201 == 3'b000;
  /* TG68KdotC_Kernel.vhd:3088:65  */
  assign n7206 = n7203 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7208 = n7225 ? 2'b01 : n1903;
  assign n7209 = {n7206, n7200};
  assign n7210 = n1785[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:3082:57  */
  assign n7211 = n7198 ? n7210 : n7209;
  assign n7212 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7213 = n7230 ? 1'b1 : n7212;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7215 = n7236 ? 7'b1001111 : n2057;
  /* TG68KdotC_Kernel.vhd:3081:49  */
  assign n7216 = n7198 & decodeopc;
  assign n7217 = n1785[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7218 = n7228 ? n7211 : n7217;
  /* TG68KdotC_Kernel.vhd:3081:49  */
  assign n7220 = n7198 & decodeopc;
  /* TG68KdotC_Kernel.vhd:3081:49  */
  assign n7221 = n7198 & decodeopc;
  /* TG68KdotC_Kernel.vhd:3097:71  */
  assign n7223 = opcode[4:3]; // extract
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7225 = n7216 & n7194;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7226 = n7194 ? n7196 : n7223;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7228 = decodeopc & n7194;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7230 = n7220 & n7194;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7232 = n7194 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7233 = n7194 ? 1'b1 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7235 = n7194 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3077:41  */
  assign n7236 = n7221 & n7194;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7237 = n7155 & n6891;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7238 = n6891 ? n7156 : n7208;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7241 = n6891 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7243 = n6891 ? n7157 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7245 = n6891 ? n7159 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7247 = n6891 ? n7161 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7249 = n6891 ? n7163 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7251 = n6891 ? n7165 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7253 = n6891 ? n7167 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7254 = n6891 ? n6913 : n7226;
  assign n7255 = n1785[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7256 = n6891 ? n7255 : n7218;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7258 = n6891 ? n7169 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7260 = n6891 ? n7170 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7262 = n6891 ? n7172 : 1'b0;
  assign n7263 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7264 = n6891 ? n7263 : n7213;
  assign n7265 = n1788[29]; // extract
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7266 = n6891 ? n7174 : n7265;
  assign n7267 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7268 = n6891 ? n7176 : n7267;
  assign n7269 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7270 = n6891 ? n7178 : n7269;
  assign n7271 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7272 = n6891 ? n7180 : n7271;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7274 = n6891 ? 1'b0 : n7232;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7276 = n6891 ? n7181 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7277 = n6891 ? n7183 : n7233;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7279 = n6891 ? n7185 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7280 = n6891 ? n7187 : n7235;
  /* TG68KdotC_Kernel.vhd:2995:33  */
  assign n7281 = n6891 ? n7188 : n7215;
  /* TG68KdotC_Kernel.vhd:2994:25  */
  assign n7283 = n2058 == 4'b1110;
  /* TG68KdotC_Kernel.vhd:3104:39  */
  assign n7284 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3104:57  */
  assign n7285 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:3104:69  */
  assign n7287 = n7285 == 3'b100;
  /* TG68KdotC_Kernel.vhd:3104:47  */
  assign n7288 = n7287 & n7284;
  /* TG68KdotC_Kernel.vhd:3105:50  */
  assign n7289 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:3105:62  */
  assign n7291 = n7289 != 2'b00;
  /* TG68KdotC_Kernel.vhd:3105:79  */
  assign n7292 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3105:91  */
  assign n7294 = n7292 != 3'b011;
  /* TG68KdotC_Kernel.vhd:3105:69  */
  assign n7295 = n7294 & n7291;
  /* TG68KdotC_Kernel.vhd:3106:51  */
  assign n7296 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3106:63  */
  assign n7298 = n7296 != 3'b111;
  /* TG68KdotC_Kernel.vhd:3106:80  */
  assign n7299 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:3106:92  */
  assign n7301 = n7299 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3106:71  */
  assign n7302 = n7298 | n7301;
  /* TG68KdotC_Kernel.vhd:3105:99  */
  assign n7303 = n7302 & n7295;
  /* TG68KdotC_Kernel.vhd:3107:58  */
  assign n7304 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3107:71  */
  assign n7306 = n7304 != 3'b000;
  /* TG68KdotC_Kernel.vhd:3109:74  */
  assign n7307 = opcode[5]; // extract
  /* TG68KdotC_Kernel.vhd:3109:77  */
  assign n7308 = ~n7307;
  /* TG68KdotC_Kernel.vhd:3109:92  */
  assign n7309 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:3109:104  */
  assign n7311 = n7309 != 2'b01;
  /* TG68KdotC_Kernel.vhd:3109:82  */
  assign n7312 = n7311 & n7308;
  /* TG68KdotC_Kernel.vhd:3109:65  */
  assign n7315 = n7312 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3109:65  */
  assign n7318 = n7312 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3108:57  */
  assign n7320 = svmode ? n7315 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3108:57  */
  assign n7323 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3108:57  */
  assign n7325 = svmode ? n7318 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3123:57  */
  assign n7328 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3123:57  */
  assign n7331 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3107:49  */
  assign n7333 = n7306 ? n7320 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3107:49  */
  assign n7334 = n7306 ? n7323 : n7328;
  /* TG68KdotC_Kernel.vhd:3107:49  */
  assign n7335 = n7306 ? n7325 : n7331;
  /* TG68KdotC_Kernel.vhd:3105:41  */
  assign n7337 = n7303 ? n7333 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3105:41  */
  assign n7339 = n7303 ? n7334 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3105:41  */
  assign n7341 = n7303 ? n7335 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3135:42  */
  assign n7342 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3135:60  */
  assign n7343 = opcode[8:6]; // extract
  /* TG68KdotC_Kernel.vhd:3135:72  */
  assign n7345 = n7343 == 3'b101;
  /* TG68KdotC_Kernel.vhd:3135:50  */
  assign n7346 = n7345 & n7342;
  /* TG68KdotC_Kernel.vhd:3136:50  */
  assign n7347 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:3136:62  */
  assign n7349 = n7347 != 2'b00;
  /* TG68KdotC_Kernel.vhd:3136:79  */
  assign n7350 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3136:91  */
  assign n7352 = n7350 != 3'b100;
  /* TG68KdotC_Kernel.vhd:3136:69  */
  assign n7353 = n7352 & n7349;
  /* TG68KdotC_Kernel.vhd:3137:51  */
  assign n7354 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3137:63  */
  assign n7356 = n7354 != 3'b111;
  /* TG68KdotC_Kernel.vhd:3137:81  */
  assign n7357 = opcode[2:1]; // extract
  /* TG68KdotC_Kernel.vhd:3137:93  */
  assign n7359 = n7357 != 2'b11;
  /* TG68KdotC_Kernel.vhd:3138:50  */
  assign n7360 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:3138:62  */
  assign n7362 = n7360 != 3'b101;
  /* TG68KdotC_Kernel.vhd:3137:100  */
  assign n7363 = n7362 & n7359;
  /* TG68KdotC_Kernel.vhd:3137:71  */
  assign n7364 = n7356 | n7363;
  /* TG68KdotC_Kernel.vhd:3136:99  */
  assign n7365 = n7364 & n7353;
  /* TG68KdotC_Kernel.vhd:3139:58  */
  assign n7366 = opcode[5:1]; // extract
  /* TG68KdotC_Kernel.vhd:3139:70  */
  assign n7368 = n7366 != 5'b11110;
  /* TG68KdotC_Kernel.vhd:3140:66  */
  assign n7369 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3140:79  */
  assign n7371 = n7369 == 3'b001;
  /* TG68KdotC_Kernel.vhd:3140:95  */
  assign n7372 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3140:108  */
  assign n7374 = n7372 == 3'b010;
  /* TG68KdotC_Kernel.vhd:3140:86  */
  assign n7375 = n7371 | n7374;
  /* TG68KdotC_Kernel.vhd:3142:82  */
  assign n7376 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3142:94  */
  assign n7378 = n7376 == 3'b101;
  /* TG68KdotC_Kernel.vhd:3142:73  */
  assign n7381 = n7378 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3142:73  */
  assign n7384 = n7378 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3141:65  */
  assign n7386 = svmode ? n7381 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3141:65  */
  assign n7389 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3141:65  */
  assign n7391 = svmode ? n7384 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3155:65  */
  assign n7394 = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3155:65  */
  assign n7397 = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3140:57  */
  assign n7399 = n7375 ? n7386 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3140:57  */
  assign n7400 = n7375 ? n7389 : n7394;
  /* TG68KdotC_Kernel.vhd:3140:57  */
  assign n7401 = n7375 ? n7391 : n7397;
  /* TG68KdotC_Kernel.vhd:3139:49  */
  assign n7403 = n7368 ? n7399 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3139:49  */
  assign n7405 = n7368 ? n7400 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3139:49  */
  assign n7407 = n7368 ? n7401 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3136:41  */
  assign n7409 = n7365 ? n7403 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3136:41  */
  assign n7411 = n7365 ? n7405 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3136:41  */
  assign n7413 = n7365 ? n7407 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3135:33  */
  assign n7415 = n7346 ? n7409 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3135:33  */
  assign n7417 = n7346 ? n7411 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3135:33  */
  assign n7419 = n7346 ? n7413 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3104:33  */
  assign n7420 = n7288 ? n7337 : n7415;
  /* TG68KdotC_Kernel.vhd:3104:33  */
  assign n7421 = n7288 ? n7339 : n7417;
  /* TG68KdotC_Kernel.vhd:3104:33  */
  assign n7422 = n7288 ? n7341 : n7419;
  /* TG68KdotC_Kernel.vhd:3103:25  */
  assign n7424 = n2058 == 4'b1111;
  assign n7425 = {n7424, n7283, n6888, n6627, n6422, n6420, n6303, n5980, n5957, n5899, n5679, n3220, n3014};
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7426 = make_berr;
      13'b0100000000000: n7426 = make_berr;
      13'b0010000000000: n7426 = make_berr;
      13'b0001000000000: n7426 = make_berr;
      13'b0000100000000: n7426 = make_berr;
      13'b0000010000000: n7426 = make_berr;
      13'b0000001000000: n7426 = make_berr;
      13'b0000000100000: n7426 = make_berr;
      13'b0000000010000: n7426 = make_berr;
      13'b0000000001000: n7426 = n5872;
      13'b0000000000100: n7426 = n5567;
      13'b0000000000010: n7426 = make_berr;
      13'b0000000000001: n7426 = make_berr;
      default: n7426 = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7428 = n1800;
      13'b0100000000000: n7428 = n6909;
      13'b0010000000000: n7428 = n6850;
      13'b0001000000000: n7428 = n6437;
      13'b0000100000000: n7428 = n1800;
      13'b0000010000000: n7428 = n6344;
      13'b0000001000000: n7428 = n6264;
      13'b0000000100000: n7428 = n5964;
      13'b0000000010000: n7428 = 2'b10;
      13'b0000000001000: n7428 = n5873;
      13'b0000000000100: n7428 = n5568;
      13'b0000000000010: n7428 = n3179;
      13'b0000000000001: n7428 = n2953;
      default: n7428 = n1800;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7429 = datatype;
      13'b0100000000000: n7429 = datatype;
      13'b0010000000000: n7429 = datatype;
      13'b0001000000000: n7429 = datatype;
      13'b0000100000000: n7429 = datatype;
      13'b0000010000000: n7429 = datatype;
      13'b0000001000000: n7429 = n6265;
      13'b0000000100000: n7429 = datatype;
      13'b0000000010000: n7429 = datatype;
      13'b0000000001000: n7429 = datatype;
      13'b0000000000100: n7429 = datatype;
      13'b0000000000010: n7429 = datatype;
      13'b0000000000001: n7429 = datatype;
      default: n7429 = datatype;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7430 = n1903;
      13'b0100000000000: n7430 = n7238;
      13'b0010000000000: n7430 = n6851;
      13'b0001000000000: n7430 = n6596;
      13'b0000100000000: n7430 = n1903;
      13'b0000010000000: n7430 = n1903;
      13'b0000001000000: n7430 = n6012;
      13'b0000000100000: n7430 = n1903;
      13'b0000000010000: n7430 = n5948;
      13'b0000000001000: n7430 = n5874;
      13'b0000000000100: n7430 = n5569;
      13'b0000000000010: n7430 = n3169;
      13'b0000000000001: n7430 = n2954;
      default: n7430 = n1903;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7431 = n2025;
      13'b0100000000000: n7431 = n2025;
      13'b0010000000000: n7431 = n2025;
      13'b0001000000000: n7431 = n2025;
      13'b0000100000000: n7431 = n2025;
      13'b0000010000000: n7431 = n2025;
      13'b0000001000000: n7431 = n2025;
      13'b0000000100000: n7431 = n2025;
      13'b0000000010000: n7431 = n2025;
      13'b0000000001000: n7431 = n2025;
      13'b0000000000100: n7431 = n5570;
      13'b0000000000010: n7431 = n2025;
      13'b0000000000001: n7431 = n2025;
      default: n7431 = n2025;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7433 = 1'b0;
      13'b0100000000000: n7433 = 1'b0;
      13'b0010000000000: n7433 = n6853;
      13'b0001000000000: n7433 = 1'b0;
      13'b0000100000000: n7433 = 1'b0;
      13'b0000010000000: n7433 = 1'b0;
      13'b0000001000000: n7433 = n6268;
      13'b0000000100000: n7433 = 1'b0;
      13'b0000000010000: n7433 = 1'b0;
      13'b0000000001000: n7433 = 1'b0;
      13'b0000000000100: n7433 = 1'b0;
      13'b0000000000010: n7433 = 1'b0;
      13'b0000000000001: n7433 = 1'b0;
      default: n7433 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7435 = n2028;
      13'b0100000000000: n7435 = n2028;
      13'b0010000000000: n7435 = n2028;
      13'b0001000000000: n7435 = n2028;
      13'b0000100000000: n7435 = n2028;
      13'b0000010000000: n7435 = n2028;
      13'b0000001000000: n7435 = n2028;
      13'b0000000100000: n7435 = n2028;
      13'b0000000010000: n7435 = n2028;
      13'b0000000001000: n7435 = n2028;
      13'b0000000000100: n7435 = n5571;
      13'b0000000000010: n7435 = n3170;
      13'b0000000000001: n7435 = n2028;
      default: n7435 = n2028;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7437 = 1'b0;
      13'b0100000000000: n7437 = n7241;
      13'b0010000000000: n7437 = 1'b0;
      13'b0001000000000: n7437 = 1'b0;
      13'b0000100000000: n7437 = 1'b0;
      13'b0000010000000: n7437 = 1'b0;
      13'b0000001000000: n7437 = 1'b0;
      13'b0000000100000: n7437 = 1'b0;
      13'b0000000010000: n7437 = 1'b0;
      13'b0000000001000: n7437 = n5876;
      13'b0000000000100: n7437 = 1'b0;
      13'b0000000000010: n7437 = 1'b0;
      13'b0000000000001: n7437 = 1'b0;
      default: n7437 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7440 = 1'b0;
      13'b0100000000000: n7440 = n7243;
      13'b0010000000000: n7440 = 1'b0;
      13'b0001000000000: n7440 = 1'b0;
      13'b0000100000000: n7440 = 1'b0;
      13'b0000010000000: n7440 = 1'b0;
      13'b0000001000000: n7440 = n6270;
      13'b0000000100000: n7440 = 1'b0;
      13'b0000000010000: n7440 = 1'b0;
      13'b0000000001000: n7440 = n5877;
      13'b0000000000100: n7440 = n5573;
      13'b0000000000010: n7440 = 1'b0;
      13'b0000000000001: n7440 = n2956;
      default: n7440 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7442 = n1892;
      13'b0100000000000: n7442 = n1892;
      13'b0010000000000: n7442 = n1892;
      13'b0001000000000: n7442 = n1892;
      13'b0000100000000: n7442 = n1892;
      13'b0000010000000: n7442 = n1892;
      13'b0000001000000: n7442 = n1892;
      13'b0000000100000: n7442 = n1892;
      13'b0000000010000: n7442 = n5940;
      13'b0000000001000: n7442 = n1892;
      13'b0000000000100: n7442 = n5574;
      13'b0000000000010: n7442 = n1892;
      13'b0000000000001: n7442 = n1892;
      default: n7442 = n1892;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7444 = 1'b0;
      13'b0100000000000: n7444 = 1'b0;
      13'b0010000000000: n7444 = 1'b0;
      13'b0001000000000: n7444 = 1'b0;
      13'b0000100000000: n7444 = 1'b0;
      13'b0000010000000: n7444 = 1'b0;
      13'b0000001000000: n7444 = 1'b0;
      13'b0000000100000: n7444 = 1'b0;
      13'b0000000010000: n7444 = n5951;
      13'b0000000001000: n7444 = 1'b0;
      13'b0000000000100: n7444 = n5576;
      13'b0000000000010: n7444 = 1'b0;
      13'b0000000000001: n7444 = 1'b0;
      default: n7444 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7447 = 1'b0;
      13'b0100000000000: n7447 = 1'b0;
      13'b0010000000000: n7447 = 1'b0;
      13'b0001000000000: n7447 = 1'b0;
      13'b0000100000000: n7447 = 1'b0;
      13'b0000010000000: n7447 = 1'b0;
      13'b0000001000000: n7447 = 1'b0;
      13'b0000000100000: n7447 = 1'b0;
      13'b0000000010000: n7447 = 1'b0;
      13'b0000000001000: n7447 = 1'b0;
      13'b0000000000100: n7447 = n5578;
      13'b0000000000010: n7447 = 1'b0;
      13'b0000000000001: n7447 = 1'b0;
      default: n7447 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7450 = 1'b0;
      13'b0100000000000: n7450 = n7245;
      13'b0010000000000: n7450 = 1'b0;
      13'b0001000000000: n7450 = 1'b0;
      13'b0000100000000: n7450 = 1'b0;
      13'b0000010000000: n7450 = 1'b0;
      13'b0000001000000: n7450 = 1'b0;
      13'b0000000100000: n7450 = 1'b0;
      13'b0000000010000: n7450 = 1'b0;
      13'b0000000001000: n7450 = 1'b0;
      13'b0000000000100: n7450 = n5579;
      13'b0000000000010: n7450 = 1'b0;
      13'b0000000000001: n7450 = 1'b0;
      default: n7450 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7453 = 1'b0;
      13'b0100000000000: n7453 = 1'b0;
      13'b0010000000000: n7453 = n6855;
      13'b0001000000000: n7453 = n6598;
      13'b0000100000000: n7453 = 1'b0;
      13'b0000010000000: n7453 = n6388;
      13'b0000001000000: n7453 = 1'b0;
      13'b0000000100000: n7453 = 1'b0;
      13'b0000000010000: n7453 = 1'b0;
      13'b0000000001000: n7453 = 1'b0;
      13'b0000000000100: n7453 = n5580;
      13'b0000000000010: n7453 = n3183;
      13'b0000000000001: n7453 = 1'b0;
      default: n7453 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7456 = 1'b0;
      13'b0100000000000: n7456 = n7247;
      13'b0010000000000: n7456 = n6857;
      13'b0001000000000: n7456 = n6600;
      13'b0000100000000: n7456 = 1'b0;
      13'b0000010000000: n7456 = n6390;
      13'b0000001000000: n7456 = n6271;
      13'b0000000100000: n7456 = 1'b0;
      13'b0000000010000: n7456 = 1'b0;
      13'b0000000001000: n7456 = 1'b0;
      13'b0000000000100: n7456 = n5581;
      13'b0000000000010: n7456 = n3186;
      13'b0000000000001: n7456 = 1'b0;
      default: n7456 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7459 = 1'b0;
      13'b0100000000000: n7459 = n7249;
      13'b0010000000000: n7459 = 1'b0;
      13'b0001000000000: n7459 = 1'b0;
      13'b0000100000000: n7459 = 1'b0;
      13'b0000010000000: n7459 = 1'b0;
      13'b0000001000000: n7459 = 1'b0;
      13'b0000000100000: n7459 = 1'b0;
      13'b0000000010000: n7459 = 1'b0;
      13'b0000000001000: n7459 = 1'b0;
      13'b0000000000100: n7459 = 1'b0;
      13'b0000000000010: n7459 = 1'b0;
      13'b0000000000001: n7459 = 1'b0;
      default: n7459 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7462 = 1'b0;
      13'b0100000000000: n7462 = n7251;
      13'b0010000000000: n7462 = 1'b0;
      13'b0001000000000: n7462 = 1'b0;
      13'b0000100000000: n7462 = 1'b0;
      13'b0000010000000: n7462 = 1'b0;
      13'b0000001000000: n7462 = 1'b0;
      13'b0000000100000: n7462 = 1'b0;
      13'b0000000010000: n7462 = 1'b0;
      13'b0000000001000: n7462 = 1'b0;
      13'b0000000000100: n7462 = n5583;
      13'b0000000000010: n7462 = 1'b0;
      13'b0000000000001: n7462 = n2958;
      default: n7462 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7465 = 1'b0;
      13'b0100000000000: n7465 = 1'b0;
      13'b0010000000000: n7465 = n6859;
      13'b0001000000000: n7465 = n6602;
      13'b0000100000000: n7465 = 1'b0;
      13'b0000010000000: n7465 = n6392;
      13'b0000001000000: n7465 = 1'b0;
      13'b0000000100000: n7465 = 1'b0;
      13'b0000000010000: n7465 = 1'b0;
      13'b0000000001000: n7465 = 1'b0;
      13'b0000000000100: n7465 = n5585;
      13'b0000000000010: n7465 = n3188;
      13'b0000000000001: n7465 = 1'b0;
      default: n7465 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7468 = 1'b0;
      13'b0100000000000: n7468 = n7253;
      13'b0010000000000: n7468 = 1'b0;
      13'b0001000000000: n7468 = 1'b0;
      13'b0000100000000: n7468 = 1'b0;
      13'b0000010000000: n7468 = 1'b0;
      13'b0000001000000: n7468 = 1'b0;
      13'b0000000100000: n7468 = 1'b0;
      13'b0000000010000: n7468 = 1'b0;
      13'b0000000001000: n7468 = 1'b0;
      13'b0000000000100: n7468 = n5587;
      13'b0000000000010: n7468 = 1'b0;
      13'b0000000000001: n7468 = 1'b0;
      default: n7468 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7471 = 1'b0;
      13'b0100000000000: n7471 = 1'b0;
      13'b0010000000000: n7471 = n6860;
      13'b0001000000000: n7471 = n6604;
      13'b0000100000000: n7471 = 1'b0;
      13'b0000010000000: n7471 = n6394;
      13'b0000001000000: n7471 = n6272;
      13'b0000000100000: n7471 = n5967;
      13'b0000000010000: n7471 = 1'b0;
      13'b0000000001000: n7471 = 1'b0;
      13'b0000000000100: n7471 = n5588;
      13'b0000000000010: n7471 = n3190;
      13'b0000000000001: n7471 = n2960;
      default: n7471 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7473 = n1779;
      13'b0100000000000: n7473 = n7254;
      13'b0010000000000: n7473 = n1779;
      13'b0001000000000: n7473 = n1779;
      13'b0000100000000: n7473 = n1779;
      13'b0000010000000: n7473 = n1779;
      13'b0000001000000: n7473 = n1779;
      13'b0000000100000: n7473 = n1779;
      13'b0000000010000: n7473 = n1779;
      13'b0000000001000: n7473 = n1779;
      13'b0000000000100: n7473 = n1779;
      13'b0000000000010: n7473 = n1779;
      13'b0000000000001: n7473 = n1779;
      default: n7473 = n1779;
    endcase
  assign n7474 = n5589[3:0]; // extract
  assign n7475 = n1785[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7476 = n7475;
      13'b0100000000000: n7476 = n7256;
      13'b0010000000000: n7476 = n7475;
      13'b0001000000000: n7476 = n7475;
      13'b0000100000000: n7476 = n7475;
      13'b0000010000000: n7476 = n7475;
      13'b0000001000000: n7476 = n7475;
      13'b0000000100000: n7476 = n7475;
      13'b0000000010000: n7476 = n7475;
      13'b0000000001000: n7476 = n7475;
      13'b0000000000100: n7476 = n7474;
      13'b0000000000010: n7476 = n7475;
      13'b0000000000001: n7476 = n7475;
      default: n7476 = n7475;
    endcase
  assign n7477 = n5589[5:4]; // extract
  assign n7478 = n1785[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7479 = n7478;
      13'b0100000000000: n7479 = n7478;
      13'b0010000000000: n7479 = n7478;
      13'b0001000000000: n7479 = n7478;
      13'b0000100000000: n7479 = n7478;
      13'b0000010000000: n7479 = n7478;
      13'b0000001000000: n7479 = n7478;
      13'b0000000100000: n7479 = n7478;
      13'b0000000010000: n7479 = n7478;
      13'b0000000001000: n7479 = n7478;
      13'b0000000000100: n7479 = n7477;
      13'b0000000000010: n7479 = n7478;
      13'b0000000000001: n7479 = n7478;
      default: n7479 = n7478;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7482 = 1'b0;
      13'b0100000000000: n7482 = 1'b0;
      13'b0010000000000: n7482 = 1'b0;
      13'b0001000000000: n7482 = 1'b0;
      13'b0000100000000: n7482 = 1'b0;
      13'b0000010000000: n7482 = 1'b0;
      13'b0000001000000: n7482 = 1'b0;
      13'b0000000100000: n7482 = 1'b0;
      13'b0000000010000: n7482 = 1'b0;
      13'b0000000001000: n7482 = 1'b0;
      13'b0000000000100: n7482 = n5591;
      13'b0000000000010: n7482 = 1'b0;
      13'b0000000000001: n7482 = 1'b0;
      default: n7482 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7484 = n2031;
      13'b0100000000000: n7484 = n2031;
      13'b0010000000000: n7484 = n2031;
      13'b0001000000000: n7484 = n2031;
      13'b0000100000000: n7484 = n2031;
      13'b0000010000000: n7484 = n2031;
      13'b0000001000000: n7484 = n6273;
      13'b0000000100000: n7484 = n2031;
      13'b0000000010000: n7484 = n2031;
      13'b0000000001000: n7484 = n2031;
      13'b0000000000100: n7484 = n5592;
      13'b0000000000010: n7484 = n2031;
      13'b0000000000001: n7484 = n2961;
      default: n7484 = n2031;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7487 = n7420;
      13'b0100000000000: n7487 = n7258;
      13'b0010000000000: n7487 = n6861;
      13'b0001000000000: n7487 = n6605;
      13'b0000100000000: n7487 = 1'b0;
      13'b0000010000000: n7487 = n6397;
      13'b0000001000000: n7487 = n6274;
      13'b0000000100000: n7487 = n5970;
      13'b0000000010000: n7487 = 1'b0;
      13'b0000000001000: n7487 = n5878;
      13'b0000000000100: n7487 = n5593;
      13'b0000000000010: n7487 = n3193;
      13'b0000000000001: n7487 = n2963;
      default: n7487 = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7490 = n7421;
      13'b0100000000000: n7490 = 1'b0;
      13'b0010000000000: n7490 = 1'b0;
      13'b0001000000000: n7490 = 1'b0;
      13'b0000100000000: n7490 = 1'b0;
      13'b0000010000000: n7490 = 1'b0;
      13'b0000001000000: n7490 = 1'b0;
      13'b0000000100000: n7490 = 1'b0;
      13'b0000000010000: n7490 = 1'b0;
      13'b0000000001000: n7490 = 1'b0;
      13'b0000000000100: n7490 = n5595;
      13'b0000000000010: n7490 = 1'b0;
      13'b0000000000001: n7490 = n2965;
      default: n7490 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7494 = 1'b0;
      13'b0100000000000: n7494 = 1'b0;
      13'b0010000000000: n7494 = 1'b0;
      13'b0001000000000: n7494 = 1'b0;
      13'b0000100000000: n7494 = 1'b1;
      13'b0000010000000: n7494 = 1'b0;
      13'b0000001000000: n7494 = 1'b0;
      13'b0000000100000: n7494 = 1'b0;
      13'b0000000010000: n7494 = 1'b0;
      13'b0000000001000: n7494 = 1'b0;
      13'b0000000000100: n7494 = 1'b0;
      13'b0000000000010: n7494 = 1'b0;
      13'b0000000000001: n7494 = 1'b0;
      default: n7494 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7497 = n7422;
      13'b0100000000000: n7497 = 1'b0;
      13'b0010000000000: n7497 = 1'b0;
      13'b0001000000000: n7497 = 1'b0;
      13'b0000100000000: n7497 = 1'b0;
      13'b0000010000000: n7497 = 1'b0;
      13'b0000001000000: n7497 = 1'b0;
      13'b0000000100000: n7497 = 1'b0;
      13'b0000000010000: n7497 = 1'b0;
      13'b0000000001000: n7497 = 1'b0;
      13'b0000000000100: n7497 = 1'b0;
      13'b0000000000010: n7497 = 1'b0;
      13'b0000000000001: n7497 = 1'b0;
      default: n7497 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7500 = 1'b0;
      13'b0100000000000: n7500 = 1'b0;
      13'b0010000000000: n7500 = 1'b0;
      13'b0001000000000: n7500 = 1'b0;
      13'b0000100000000: n7500 = 1'b0;
      13'b0000010000000: n7500 = 1'b0;
      13'b0000001000000: n7500 = 1'b0;
      13'b0000000100000: n7500 = 1'b0;
      13'b0000000010000: n7500 = 1'b0;
      13'b0000000001000: n7500 = 1'b0;
      13'b0000000000100: n7500 = n5597;
      13'b0000000000010: n7500 = 1'b0;
      13'b0000000000001: n7500 = 1'b0;
      default: n7500 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7503 = 1'b0;
      13'b0100000000000: n7503 = 1'b0;
      13'b0010000000000: n7503 = 1'b0;
      13'b0001000000000: n7503 = 1'b0;
      13'b0000100000000: n7503 = 1'b0;
      13'b0000010000000: n7503 = 1'b0;
      13'b0000001000000: n7503 = 1'b0;
      13'b0000000100000: n7503 = 1'b0;
      13'b0000000010000: n7503 = 1'b0;
      13'b0000000001000: n7503 = n5880;
      13'b0000000000100: n7503 = n5599;
      13'b0000000000010: n7503 = 1'b0;
      13'b0000000000001: n7503 = 1'b0;
      default: n7503 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7509 = 1'b1;
      13'b0100000000000: n7509 = n7260;
      13'b0010000000000: n7509 = n6862;
      13'b0001000000000: n7509 = n6606;
      13'b0000100000000: n7509 = 1'b1;
      13'b0000010000000: n7509 = n6400;
      13'b0000001000000: n7509 = n6275;
      13'b0000000100000: n7509 = n5973;
      13'b0000000010000: n7509 = 1'b0;
      13'b0000000001000: n7509 = n5881;
      13'b0000000000100: n7509 = n5600;
      13'b0000000000010: n7509 = n3196;
      13'b0000000000001: n7509 = n2967;
      default: n7509 = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7512 = 1'b0;
      13'b0100000000000: n7512 = 1'b0;
      13'b0010000000000: n7512 = 1'b0;
      13'b0001000000000: n7512 = 1'b0;
      13'b0000100000000: n7512 = 1'b0;
      13'b0000010000000: n7512 = 1'b0;
      13'b0000001000000: n7512 = 1'b0;
      13'b0000000100000: n7512 = 1'b0;
      13'b0000000010000: n7512 = 1'b0;
      13'b0000000001000: n7512 = 1'b0;
      13'b0000000000100: n7512 = n5602;
      13'b0000000000010: n7512 = 1'b0;
      13'b0000000000001: n7512 = 1'b0;
      default: n7512 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7515 = 1'b0;
      13'b0100000000000: n7515 = n7262;
      13'b0010000000000: n7515 = n6864;
      13'b0001000000000: n7515 = n6607;
      13'b0000100000000: n7515 = 1'b0;
      13'b0000010000000: n7515 = n6403;
      13'b0000001000000: n7515 = n6277;
      13'b0000000100000: n7515 = 1'b0;
      13'b0000000010000: n7515 = 1'b0;
      13'b0000000001000: n7515 = n5882;
      13'b0000000000100: n7515 = n5603;
      13'b0000000000010: n7515 = n3199;
      13'b0000000000001: n7515 = n2969;
      default: n7515 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7518 = 1'b0;
      13'b0100000000000: n7518 = 1'b0;
      13'b0010000000000: n7518 = n6866;
      13'b0001000000000: n7518 = n6609;
      13'b0000100000000: n7518 = 1'b0;
      13'b0000010000000: n7518 = n6405;
      13'b0000001000000: n7518 = n6279;
      13'b0000000100000: n7518 = 1'b0;
      13'b0000000010000: n7518 = 1'b0;
      13'b0000000001000: n7518 = 1'b0;
      13'b0000000000100: n7518 = 1'b0;
      13'b0000000000010: n7518 = 1'b0;
      13'b0000000000001: n7518 = 1'b0;
      default: n7518 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7521 = 1'b0;
      13'b0100000000000: n7521 = 1'b0;
      13'b0010000000000: n7521 = n6868;
      13'b0001000000000: n7521 = 1'b0;
      13'b0000100000000: n7521 = 1'b0;
      13'b0000010000000: n7521 = n6407;
      13'b0000001000000: n7521 = n6281;
      13'b0000000100000: n7521 = 1'b0;
      13'b0000000010000: n7521 = 1'b0;
      13'b0000000001000: n7521 = 1'b0;
      13'b0000000000100: n7521 = 1'b0;
      13'b0000000000010: n7521 = 1'b0;
      13'b0000000000001: n7521 = 1'b0;
      default: n7521 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7524 = 1'b0;
      13'b0100000000000: n7524 = 1'b0;
      13'b0010000000000: n7524 = 1'b0;
      13'b0001000000000: n7524 = 1'b0;
      13'b0000100000000: n7524 = 1'b0;
      13'b0000010000000: n7524 = 1'b0;
      13'b0000001000000: n7524 = 1'b0;
      13'b0000000100000: n7524 = 1'b0;
      13'b0000000010000: n7524 = 1'b0;
      13'b0000000001000: n7524 = 1'b0;
      13'b0000000000100: n7524 = 1'b0;
      13'b0000000000010: n7524 = 1'b0;
      13'b0000000000001: n7524 = n2971;
      default: n7524 = 1'b0;
    endcase
  assign n7526 = n1788[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7527 = n7526;
      13'b0100000000000: n7527 = n7526;
      13'b0010000000000: n7527 = n7526;
      13'b0001000000000: n7527 = n7526;
      13'b0000100000000: n7527 = n7526;
      13'b0000010000000: n7527 = n7526;
      13'b0000001000000: n7527 = n7526;
      13'b0000000100000: n7527 = n7526;
      13'b0000000010000: n7527 = n7526;
      13'b0000000001000: n7527 = n7526;
      13'b0000000000100: n7527 = n5609;
      13'b0000000000010: n7527 = n7526;
      13'b0000000000001: n7527 = n7526;
      default: n7527 = n7526;
    endcase
  assign n7528 = n1788[19:17]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7529 = n7528;
      13'b0100000000000: n7529 = n7528;
      13'b0010000000000: n7529 = n7528;
      13'b0001000000000: n7529 = n7528;
      13'b0000100000000: n7529 = n7528;
      13'b0000010000000: n7529 = n7528;
      13'b0000001000000: n7529 = n7528;
      13'b0000000100000: n7529 = n7528;
      13'b0000000010000: n7529 = n7528;
      13'b0000000001000: n7529 = n7528;
      13'b0000000000100: n7529 = n7528;
      13'b0000000000010: n7529 = n7528;
      13'b0000000000001: n7529 = n2975;
      default: n7529 = n7528;
    endcase
  assign n7530 = n1788[20]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7531 = n7530;
      13'b0100000000000: n7531 = n7530;
      13'b0010000000000: n7531 = n7530;
      13'b0001000000000: n7531 = n7530;
      13'b0000100000000: n7531 = n7530;
      13'b0000010000000: n7531 = n7530;
      13'b0000001000000: n7531 = n7530;
      13'b0000000100000: n7531 = n7530;
      13'b0000000010000: n7531 = n7530;
      13'b0000000001000: n7531 = n7530;
      13'b0000000000100: n7531 = n5611;
      13'b0000000000010: n7531 = n7530;
      13'b0000000000001: n7531 = n7530;
      default: n7531 = n7530;
    endcase
  assign n7532 = n1788[24]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7533 = n7532;
      13'b0100000000000: n7533 = n7264;
      13'b0010000000000: n7533 = n7532;
      13'b0001000000000: n7533 = n7532;
      13'b0000100000000: n7533 = n7532;
      13'b0000010000000: n7533 = n7532;
      13'b0000001000000: n7533 = n7532;
      13'b0000000100000: n7533 = n7532;
      13'b0000000010000: n7533 = n7532;
      13'b0000000001000: n7533 = n7532;
      13'b0000000000100: n7533 = n5613;
      13'b0000000000010: n7533 = n7532;
      13'b0000000000001: n7533 = n7532;
      default: n7533 = n7532;
    endcase
  assign n7534 = n1788[26]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7535 = n7534;
      13'b0100000000000: n7535 = n7534;
      13'b0010000000000: n7535 = n7534;
      13'b0001000000000: n7535 = n7534;
      13'b0000100000000: n7535 = n7534;
      13'b0000010000000: n7535 = n7534;
      13'b0000001000000: n7535 = n7534;
      13'b0000000100000: n7535 = n7534;
      13'b0000000010000: n7535 = n7534;
      13'b0000000001000: n7535 = n7534;
      13'b0000000000100: n7535 = n7534;
      13'b0000000000010: n7535 = n7534;
      13'b0000000000001: n7535 = n2977;
      default: n7535 = n7534;
    endcase
  assign n7536 = n1788[29]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7537 = n7536;
      13'b0100000000000: n7537 = n7266;
      13'b0010000000000: n7537 = n7536;
      13'b0001000000000: n7537 = n7536;
      13'b0000100000000: n7537 = n7536;
      13'b0000010000000: n7537 = n7536;
      13'b0000001000000: n7537 = n7536;
      13'b0000000100000: n7537 = n7536;
      13'b0000000010000: n7537 = n7536;
      13'b0000000001000: n7537 = n7536;
      13'b0000000000100: n7537 = n7536;
      13'b0000000000010: n7537 = n7536;
      13'b0000000000001: n7537 = n7536;
      default: n7537 = n7536;
    endcase
  assign n7538 = n1788[34]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7539 = n7538;
      13'b0100000000000: n7539 = n7538;
      13'b0010000000000: n7539 = n6870;
      13'b0001000000000: n7539 = n7538;
      13'b0000100000000: n7539 = n7538;
      13'b0000010000000: n7539 = n7538;
      13'b0000001000000: n7539 = n7538;
      13'b0000000100000: n7539 = n7538;
      13'b0000000010000: n7539 = n7538;
      13'b0000000001000: n7539 = n7538;
      13'b0000000000100: n7539 = n5615;
      13'b0000000000010: n7539 = n7538;
      13'b0000000000001: n7539 = n7538;
      default: n7539 = n7538;
    endcase
  assign n7540 = n1788[36]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7541 = n7540;
      13'b0100000000000: n7541 = n7540;
      13'b0010000000000: n7541 = n7540;
      13'b0001000000000: n7541 = n7540;
      13'b0000100000000: n7541 = n7540;
      13'b0000010000000: n7541 = n7540;
      13'b0000001000000: n7541 = n7540;
      13'b0000000100000: n7541 = n7540;
      13'b0000000010000: n7541 = n7540;
      13'b0000000001000: n7541 = n7540;
      13'b0000000000100: n7541 = n5617;
      13'b0000000000010: n7541 = n7540;
      13'b0000000000001: n7541 = n7540;
      default: n7541 = n7540;
    endcase
  assign n7542 = n1788[37]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7543 = n7542;
      13'b0100000000000: n7543 = n7542;
      13'b0010000000000: n7543 = n7542;
      13'b0001000000000: n7543 = n7542;
      13'b0000100000000: n7543 = n7542;
      13'b0000010000000: n7543 = n7542;
      13'b0000001000000: n7543 = n7542;
      13'b0000000100000: n7543 = n7542;
      13'b0000000010000: n7543 = n7542;
      13'b0000000001000: n7543 = n7542;
      13'b0000000000100: n7543 = n7542;
      13'b0000000000010: n7543 = n7542;
      13'b0000000000001: n7543 = n2979;
      default: n7543 = n7542;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7544 = n1884;
      13'b0100000000000: n7544 = n1884;
      13'b0010000000000: n7544 = n1884;
      13'b0001000000000: n7544 = n6610;
      13'b0000100000000: n7544 = n1884;
      13'b0000010000000: n7544 = n1884;
      13'b0000001000000: n7544 = n1884;
      13'b0000000100000: n7544 = n1884;
      13'b0000000010000: n7544 = n1884;
      13'b0000000001000: n7544 = n1884;
      13'b0000000000100: n7544 = n1884;
      13'b0000000000010: n7544 = n1884;
      13'b0000000000001: n7544 = n1884;
      default: n7544 = n1884;
    endcase
  assign n7545 = n1788[39]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7546 = n7545;
      13'b0100000000000: n7546 = n7545;
      13'b0010000000000: n7546 = n7545;
      13'b0001000000000: n7546 = n7545;
      13'b0000100000000: n7546 = n7545;
      13'b0000010000000: n7546 = n7545;
      13'b0000001000000: n7546 = n7545;
      13'b0000000100000: n7546 = n7545;
      13'b0000000010000: n7546 = n7545;
      13'b0000000001000: n7546 = n7545;
      13'b0000000000100: n7546 = n7545;
      13'b0000000000010: n7546 = n7545;
      13'b0000000000001: n7546 = n2981;
      default: n7546 = n7545;
    endcase
  assign n7547 = n1788[40]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7548 = n7547;
      13'b0100000000000: n7548 = n7547;
      13'b0010000000000: n7548 = n7547;
      13'b0001000000000: n7548 = n7547;
      13'b0000100000000: n7548 = n7547;
      13'b0000010000000: n7548 = n7547;
      13'b0000001000000: n7548 = n7547;
      13'b0000000100000: n7548 = n7547;
      13'b0000000010000: n7548 = n7547;
      13'b0000000001000: n7548 = n7547;
      13'b0000000000100: n7548 = n5619;
      13'b0000000000010: n7548 = n3173;
      13'b0000000000001: n7548 = n7547;
      default: n7548 = n7547;
    endcase
  assign n7549 = n2983[0]; // extract
  assign n7550 = n1788[42]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7551 = n7550;
      13'b0100000000000: n7551 = n7268;
      13'b0010000000000: n7551 = n7550;
      13'b0001000000000: n7551 = n7550;
      13'b0000100000000: n7551 = n7550;
      13'b0000010000000: n7551 = n7550;
      13'b0000001000000: n7551 = n7550;
      13'b0000000100000: n7551 = n7550;
      13'b0000000010000: n7551 = n7550;
      13'b0000000001000: n7551 = n7550;
      13'b0000000000100: n7551 = n5621;
      13'b0000000000010: n7551 = n7550;
      13'b0000000000001: n7551 = n7549;
      default: n7551 = n7550;
    endcase
  assign n7552 = n2983[1]; // extract
  assign n7553 = n1788[43]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7554 = n7553;
      13'b0100000000000: n7554 = n7553;
      13'b0010000000000: n7554 = n7553;
      13'b0001000000000: n7554 = n7553;
      13'b0000100000000: n7554 = n7553;
      13'b0000010000000: n7554 = n7553;
      13'b0000001000000: n7554 = n7553;
      13'b0000000100000: n7554 = n7553;
      13'b0000000010000: n7554 = n7553;
      13'b0000000001000: n7554 = n7553;
      13'b0000000000100: n7554 = n5623;
      13'b0000000000010: n7554 = n7553;
      13'b0000000000001: n7554 = n7552;
      default: n7554 = n7553;
    endcase
  assign n7555 = n1788[44]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7556 = n7555;
      13'b0100000000000: n7556 = n7555;
      13'b0010000000000: n7556 = n7555;
      13'b0001000000000: n7556 = n7555;
      13'b0000100000000: n7556 = n7555;
      13'b0000010000000: n7556 = n7555;
      13'b0000001000000: n7556 = n6283;
      13'b0000000100000: n7556 = n7555;
      13'b0000000010000: n7556 = n7555;
      13'b0000000001000: n7556 = n7555;
      13'b0000000000100: n7556 = n5625;
      13'b0000000000010: n7556 = n7555;
      13'b0000000000001: n7556 = n7555;
      default: n7556 = n7555;
    endcase
  assign n7557 = n3174[0]; // extract
  assign n7558 = n5629[0]; // extract
  assign n7559 = n2043[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7560 = n7559;
      13'b0100000000000: n7560 = n7559;
      13'b0010000000000: n7560 = n7559;
      13'b0001000000000: n7560 = n6612;
      13'b0000100000000: n7560 = n7559;
      13'b0000010000000: n7560 = n7559;
      13'b0000001000000: n7560 = n7559;
      13'b0000000100000: n7560 = n7559;
      13'b0000000010000: n7560 = n7559;
      13'b0000000001000: n7560 = n7559;
      13'b0000000000100: n7560 = n7558;
      13'b0000000000010: n7560 = n7557;
      13'b0000000000001: n7560 = n7559;
      default: n7560 = n7559;
    endcase
  assign n7561 = n3174[1]; // extract
  assign n7562 = n5629[1]; // extract
  assign n7563 = n2043[1]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7564 = n7563;
      13'b0100000000000: n7564 = n7563;
      13'b0010000000000: n7564 = n7563;
      13'b0001000000000: n7564 = n7563;
      13'b0000100000000: n7564 = n7563;
      13'b0000010000000: n7564 = n7563;
      13'b0000001000000: n7564 = n7563;
      13'b0000000100000: n7564 = n7563;
      13'b0000000010000: n7564 = n5944;
      13'b0000000001000: n7564 = n7563;
      13'b0000000000100: n7564 = n7562;
      13'b0000000000010: n7564 = n7561;
      13'b0000000000001: n7564 = n7563;
      default: n7564 = n7563;
    endcase
  assign n7565 = n5629[2]; // extract
  assign n7566 = n1788[48]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7567 = n7566;
      13'b0100000000000: n7567 = n7566;
      13'b0010000000000: n7567 = n7566;
      13'b0001000000000: n7567 = n7566;
      13'b0000100000000: n7567 = n7566;
      13'b0000010000000: n7567 = n7566;
      13'b0000001000000: n7567 = n7566;
      13'b0000000100000: n7567 = n7566;
      13'b0000000010000: n7567 = n7566;
      13'b0000000001000: n7567 = n7566;
      13'b0000000000100: n7567 = n7565;
      13'b0000000000010: n7567 = n7566;
      13'b0000000000001: n7567 = n7566;
      default: n7567 = n7566;
    endcase
  assign n7568 = n3206[0]; // extract
  assign n7569 = n1788[49]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7570 = n7569;
      13'b0100000000000: n7570 = n7569;
      13'b0010000000000: n7570 = n7569;
      13'b0001000000000: n7570 = n7569;
      13'b0000100000000: n7570 = n7569;
      13'b0000010000000: n7570 = n6383;
      13'b0000001000000: n7570 = n6285;
      13'b0000000100000: n7570 = n7569;
      13'b0000000010000: n7570 = n7569;
      13'b0000000001000: n7570 = n5884;
      13'b0000000000100: n7570 = n5631;
      13'b0000000000010: n7570 = n7568;
      13'b0000000000001: n7570 = n2985;
      default: n7570 = n7569;
    endcase
  assign n7571 = n3206[1]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7572 = n2045;
      13'b0100000000000: n7572 = n2045;
      13'b0010000000000: n7572 = n2045;
      13'b0001000000000: n7572 = n6613;
      13'b0000100000000: n7572 = n2045;
      13'b0000010000000: n7572 = n2045;
      13'b0000001000000: n7572 = n2045;
      13'b0000000100000: n7572 = n2045;
      13'b0000000010000: n7572 = n2045;
      13'b0000000001000: n7572 = n2045;
      13'b0000000000100: n7572 = n2045;
      13'b0000000000010: n7572 = n7571;
      13'b0000000000001: n7572 = n2987;
      default: n7572 = n2045;
    endcase
  assign n7573 = n5634[1:0]; // extract
  assign n7574 = n1788[52:51]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7575 = n7574;
      13'b0100000000000: n7575 = n7574;
      13'b0010000000000: n7575 = n7574;
      13'b0001000000000: n7575 = n7574;
      13'b0000100000000: n7575 = n7574;
      13'b0000010000000: n7575 = n7574;
      13'b0000001000000: n7575 = n7574;
      13'b0000000100000: n7575 = n7574;
      13'b0000000010000: n7575 = n7574;
      13'b0000000001000: n7575 = n7574;
      13'b0000000000100: n7575 = n7573;
      13'b0000000000010: n7575 = n7574;
      13'b0000000000001: n7575 = n2989;
      default: n7575 = n7574;
    endcase
  assign n7576 = n5634[2]; // extract
  assign n7577 = n1788[53]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7578 = n7577;
      13'b0100000000000: n7578 = n7577;
      13'b0010000000000: n7578 = n7577;
      13'b0001000000000: n7578 = n7577;
      13'b0000100000000: n7578 = n7577;
      13'b0000010000000: n7578 = n7577;
      13'b0000001000000: n7578 = n7577;
      13'b0000000100000: n7578 = n7577;
      13'b0000000010000: n7578 = n7577;
      13'b0000000001000: n7578 = n5691;
      13'b0000000000100: n7578 = n7576;
      13'b0000000000010: n7578 = n7577;
      13'b0000000000001: n7578 = n7577;
      default: n7578 = n7577;
    endcase
  assign n7579 = n5634[3]; // extract
  assign n7580 = n1788[54]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7581 = n7580;
      13'b0100000000000: n7581 = n7580;
      13'b0010000000000: n7581 = n7580;
      13'b0001000000000: n7581 = n7580;
      13'b0000100000000: n7581 = n7580;
      13'b0000010000000: n7581 = n7580;
      13'b0000001000000: n7581 = n7580;
      13'b0000000100000: n7581 = n7580;
      13'b0000000010000: n7581 = n7580;
      13'b0000000001000: n7581 = n7580;
      13'b0000000000100: n7581 = n7579;
      13'b0000000000010: n7581 = n7580;
      13'b0000000000001: n7581 = n7580;
      default: n7581 = n7580;
    endcase
  assign n7582 = n2991[0]; // extract
  assign n7583 = n5634[4]; // extract
  assign n7584 = n1788[55]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7585 = n7584;
      13'b0100000000000: n7585 = n7270;
      13'b0010000000000: n7585 = n7584;
      13'b0001000000000: n7585 = n7584;
      13'b0000100000000: n7585 = n7584;
      13'b0000010000000: n7585 = n7584;
      13'b0000001000000: n7585 = n7584;
      13'b0000000100000: n7585 = n7584;
      13'b0000000010000: n7585 = n7584;
      13'b0000000001000: n7585 = n7584;
      13'b0000000000100: n7585 = n7583;
      13'b0000000000010: n7585 = n7584;
      13'b0000000000001: n7585 = n7582;
      default: n7585 = n7584;
    endcase
  assign n7586 = n2991[1]; // extract
  assign n7587 = n1788[56]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7588 = n7587;
      13'b0100000000000: n7588 = n7587;
      13'b0010000000000: n7588 = n7587;
      13'b0001000000000: n7588 = n6614;
      13'b0000100000000: n7588 = n7587;
      13'b0000010000000: n7588 = n6337;
      13'b0000001000000: n7588 = n6287;
      13'b0000000100000: n7588 = n7587;
      13'b0000000010000: n7588 = n7587;
      13'b0000000001000: n7588 = n5888;
      13'b0000000000100: n7588 = n5636;
      13'b0000000000010: n7588 = n7587;
      13'b0000000000001: n7588 = n7586;
      default: n7588 = n7587;
    endcase
  assign n7589 = n1788[60:57]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7590 = n7589;
      13'b0100000000000: n7590 = n7589;
      13'b0010000000000: n7590 = n7589;
      13'b0001000000000: n7590 = n7589;
      13'b0000100000000: n7590 = n7589;
      13'b0000010000000: n7590 = n7589;
      13'b0000001000000: n7590 = n7589;
      13'b0000000100000: n7590 = n7589;
      13'b0000000010000: n7590 = n7589;
      13'b0000000001000: n7590 = n7589;
      13'b0000000000100: n7590 = n5639;
      13'b0000000000010: n7590 = n7589;
      13'b0000000000001: n7590 = n7589;
      default: n7590 = n7589;
    endcase
  assign n7591 = n1788[61]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7592 = n7591;
      13'b0100000000000: n7592 = n7591;
      13'b0010000000000: n7592 = n6872;
      13'b0001000000000: n7592 = n7591;
      13'b0000100000000: n7592 = n7591;
      13'b0000010000000: n7592 = n7591;
      13'b0000001000000: n7592 = n7591;
      13'b0000000100000: n7592 = n7591;
      13'b0000000010000: n7592 = n7591;
      13'b0000000001000: n7592 = n7591;
      13'b0000000000100: n7592 = n7591;
      13'b0000000000010: n7592 = n7591;
      13'b0000000000001: n7592 = n7591;
      default: n7592 = n7591;
    endcase
  assign n7593 = n1788[67]; // extract
  assign n7594 = {n7593, n1896, n2055};
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7595 = n7594;
      13'b0100000000000: n7595 = n7594;
      13'b0010000000000: n7595 = n7594;
      13'b0001000000000: n7595 = n7594;
      13'b0000100000000: n7595 = n7594;
      13'b0000010000000: n7595 = n7594;
      13'b0000001000000: n7595 = n7594;
      13'b0000000100000: n7595 = n7594;
      13'b0000000010000: n7595 = n7594;
      13'b0000000001000: n7595 = n7594;
      13'b0000000000100: n7595 = n5642;
      13'b0000000000010: n7595 = n7594;
      13'b0000000000001: n7595 = n7594;
      default: n7595 = n7594;
    endcase
  assign n7596 = n1788[69]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7597 = n7596;
      13'b0100000000000: n7597 = n7596;
      13'b0010000000000: n7597 = n7596;
      13'b0001000000000: n7597 = n7596;
      13'b0000100000000: n7597 = n7596;
      13'b0000010000000: n7597 = n7596;
      13'b0000001000000: n7597 = n7596;
      13'b0000000100000: n7597 = n7596;
      13'b0000000010000: n7597 = n7596;
      13'b0000000001000: n7597 = n7596;
      13'b0000000000100: n7597 = n5644;
      13'b0000000000010: n7597 = n7596;
      13'b0000000000001: n7597 = n7596;
      default: n7597 = n7596;
    endcase
  assign n7598 = n1788[71]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7599 = n7598;
      13'b0100000000000: n7599 = n7272;
      13'b0010000000000: n7599 = n7598;
      13'b0001000000000: n7599 = n7598;
      13'b0000100000000: n7599 = n7598;
      13'b0000010000000: n7599 = n7598;
      13'b0000001000000: n7599 = n7598;
      13'b0000000100000: n7599 = n7598;
      13'b0000000010000: n7599 = n7598;
      13'b0000000001000: n7599 = n7598;
      13'b0000000000100: n7599 = n5646;
      13'b0000000000010: n7599 = n7598;
      13'b0000000000001: n7599 = n2993;
      default: n7599 = n7598;
    endcase
  assign n7600 = n5649[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7601 = n2048;
      13'b0100000000000: n7601 = n2048;
      13'b0010000000000: n7601 = n2048;
      13'b0001000000000: n7601 = n2048;
      13'b0000100000000: n7601 = n2048;
      13'b0000010000000: n7601 = n2048;
      13'b0000001000000: n7601 = n2048;
      13'b0000000100000: n7601 = n2048;
      13'b0000000010000: n7601 = n5954;
      13'b0000000001000: n7601 = n5889;
      13'b0000000000100: n7601 = n7600;
      13'b0000000000010: n7601 = n3176;
      13'b0000000000001: n7601 = n2994;
      default: n7601 = n2048;
    endcase
  assign n7602 = n5649[1]; // extract
  assign n7603 = n1788[74]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7604 = n7603;
      13'b0100000000000: n7604 = n7603;
      13'b0010000000000: n7604 = n7603;
      13'b0001000000000: n7604 = n7603;
      13'b0000100000000: n7604 = n7603;
      13'b0000010000000: n7604 = n7603;
      13'b0000001000000: n7604 = n7603;
      13'b0000000100000: n7604 = n7603;
      13'b0000000010000: n7604 = n7603;
      13'b0000000001000: n7604 = n7603;
      13'b0000000000100: n7604 = n7602;
      13'b0000000000010: n7604 = n7603;
      13'b0000000000001: n7604 = n7603;
      default: n7604 = n7603;
    endcase
  assign n7605 = n1788[80]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7606 = n7605;
      13'b0100000000000: n7606 = n7605;
      13'b0010000000000: n7606 = n7605;
      13'b0001000000000: n7606 = n7605;
      13'b0000100000000: n7606 = n7605;
      13'b0000010000000: n7606 = n7605;
      13'b0000001000000: n7606 = n6289;
      13'b0000000100000: n7606 = n7605;
      13'b0000000010000: n7606 = n7605;
      13'b0000000001000: n7606 = n7605;
      13'b0000000000100: n7606 = n7605;
      13'b0000000000010: n7606 = n7605;
      13'b0000000000001: n7606 = n7605;
      default: n7606 = n7605;
    endcase
  assign n7607 = n1788[82]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7608 = n7607;
      13'b0100000000000: n7608 = n7607;
      13'b0010000000000: n7608 = n7607;
      13'b0001000000000: n7608 = n7607;
      13'b0000100000000: n7608 = n7607;
      13'b0000010000000: n7608 = n7607;
      13'b0000001000000: n7608 = n7607;
      13'b0000000100000: n7608 = n7607;
      13'b0000000010000: n7608 = n7607;
      13'b0000000001000: n7608 = n7607;
      13'b0000000000100: n7608 = n7607;
      13'b0000000000010: n7608 = n7607;
      13'b0000000000001: n7608 = n2996;
      default: n7608 = n7607;
    endcase
  assign n7609 = n1788[84]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7610 = n7609;
      13'b0100000000000: n7610 = n7609;
      13'b0010000000000: n7610 = n7609;
      13'b0001000000000: n7610 = n7609;
      13'b0000100000000: n7610 = n7609;
      13'b0000010000000: n7610 = n7609;
      13'b0000001000000: n7610 = n7609;
      13'b0000000100000: n7610 = n7609;
      13'b0000000010000: n7610 = n7609;
      13'b0000000001000: n7610 = n7609;
      13'b0000000000100: n7610 = n7609;
      13'b0000000000010: n7610 = n7609;
      13'b0000000000001: n7610 = n2998;
      default: n7610 = n7609;
    endcase
  assign n7611 = n1788[85]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7612 = n7611;
      13'b0100000000000: n7612 = n7611;
      13'b0010000000000: n7612 = n6874;
      13'b0001000000000: n7612 = n7611;
      13'b0000100000000: n7612 = n7611;
      13'b0000010000000: n7612 = n7611;
      13'b0000001000000: n7612 = n7611;
      13'b0000000100000: n7612 = n7611;
      13'b0000000010000: n7612 = n7611;
      13'b0000000001000: n7612 = n7611;
      13'b0000000000100: n7612 = n7611;
      13'b0000000000010: n7612 = n7611;
      13'b0000000000001: n7612 = n7611;
      default: n7612 = n7611;
    endcase
  assign n7613 = n1788[86]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7614 = n7613;
      13'b0100000000000: n7614 = n7613;
      13'b0010000000000: n7614 = n7613;
      13'b0001000000000: n7614 = n7613;
      13'b0000100000000: n7614 = n7613;
      13'b0000010000000: n7614 = n7613;
      13'b0000001000000: n7614 = n7613;
      13'b0000000100000: n7614 = n7613;
      13'b0000000010000: n7614 = n7613;
      13'b0000000001000: n7614 = n7613;
      13'b0000000000100: n7614 = n7613;
      13'b0000000000010: n7614 = n7613;
      13'b0000000000001: n7614 = n3000;
      default: n7614 = n7613;
    endcase
  assign n7617 = n1788[16:1]; // extract
  assign n7618 = n1788[21]; // extract
  assign n7619 = n1788[23]; // extract
  assign n7624 = n1788[33:30]; // extract
  assign n7626 = n1788[35]; // extract
  assign n7630 = n1788[45]; // extract
  assign n7641 = n1788[68]; // extract
  assign n7642 = n1788[72]; // extract
  assign n7643 = n1788[70]; // extract
  assign n7647 = n1788[81]; // extract
  assign n7651 = n5976[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7653 = 1'b0;
      13'b0100000000000: n7653 = 1'b0;
      13'b0010000000000: n7653 = 1'b0;
      13'b0001000000000: n7653 = 1'b0;
      13'b0000100000000: n7653 = 1'b0;
      13'b0000010000000: n7653 = 1'b0;
      13'b0000001000000: n7653 = 1'b0;
      13'b0000000100000: n7653 = n7651;
      13'b0000000010000: n7653 = 1'b0;
      13'b0000000001000: n7653 = 1'b0;
      13'b0000000000100: n7653 = n5653;
      13'b0000000000010: n7653 = n3209;
      13'b0000000000001: n7653 = n3002;
      default: n7653 = 1'b0;
    endcase
  assign n7654 = n5976[1]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7656 = 1'b0;
      13'b0100000000000: n7656 = 1'b0;
      13'b0010000000000: n7656 = 1'b0;
      13'b0001000000000: n7656 = 1'b0;
      13'b0000100000000: n7656 = 1'b0;
      13'b0000010000000: n7656 = 1'b0;
      13'b0000001000000: n7656 = 1'b0;
      13'b0000000100000: n7656 = n7654;
      13'b0000000010000: n7656 = 1'b0;
      13'b0000000001000: n7656 = 1'b0;
      13'b0000000000100: n7656 = 1'b0;
      13'b0000000000010: n7656 = 1'b0;
      13'b0000000000001: n7656 = 1'b0;
      default: n7656 = 1'b0;
    endcase
  assign n7657 = n5655[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7659 = 1'b0;
      13'b0100000000000: n7659 = 1'b0;
      13'b0010000000000: n7659 = 1'b0;
      13'b0001000000000: n7659 = 1'b0;
      13'b0000100000000: n7659 = 1'b0;
      13'b0000010000000: n7659 = 1'b0;
      13'b0000001000000: n7659 = 1'b0;
      13'b0000000100000: n7659 = 1'b0;
      13'b0000000010000: n7659 = 1'b0;
      13'b0000000001000: n7659 = 1'b0;
      13'b0000000000100: n7659 = n7657;
      13'b0000000000010: n7659 = 1'b0;
      13'b0000000000001: n7659 = 1'b0;
      default: n7659 = 1'b0;
    endcase
  assign n7660 = n5655[1]; // extract
  assign n7661 = n5891[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7663 = 1'b0;
      13'b0100000000000: n7663 = 1'b0;
      13'b0010000000000: n7663 = n6876;
      13'b0001000000000: n7663 = 1'b0;
      13'b0000100000000: n7663 = 1'b0;
      13'b0000010000000: n7663 = n6413;
      13'b0000001000000: n7663 = n6291;
      13'b0000000100000: n7663 = 1'b0;
      13'b0000000010000: n7663 = 1'b0;
      13'b0000000001000: n7663 = n7661;
      13'b0000000000100: n7663 = n7660;
      13'b0000000000010: n7663 = 1'b0;
      13'b0000000000001: n7663 = n3004;
      default: n7663 = 1'b0;
    endcase
  assign n7664 = n5891[1]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7666 = 1'b0;
      13'b0100000000000: n7666 = 1'b0;
      13'b0010000000000: n7666 = 1'b0;
      13'b0001000000000: n7666 = 1'b0;
      13'b0000100000000: n7666 = 1'b0;
      13'b0000010000000: n7666 = 1'b0;
      13'b0000001000000: n7666 = 1'b0;
      13'b0000000100000: n7666 = 1'b0;
      13'b0000000010000: n7666 = 1'b0;
      13'b0000000001000: n7666 = n7664;
      13'b0000000000100: n7666 = 1'b0;
      13'b0000000000010: n7666 = 1'b0;
      13'b0000000000001: n7666 = 1'b0;
      default: n7666 = 1'b0;
    endcase
  assign n7667 = n3006[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7669 = 1'b0;
      13'b0100000000000: n7669 = 1'b0;
      13'b0010000000000: n7669 = 1'b0;
      13'b0001000000000: n7669 = 1'b0;
      13'b0000100000000: n7669 = 1'b0;
      13'b0000010000000: n7669 = 1'b0;
      13'b0000001000000: n7669 = n6293;
      13'b0000000100000: n7669 = 1'b0;
      13'b0000000010000: n7669 = 1'b0;
      13'b0000000001000: n7669 = 1'b0;
      13'b0000000000100: n7669 = 1'b0;
      13'b0000000000010: n7669 = 1'b0;
      13'b0000000000001: n7669 = n7667;
      default: n7669 = 1'b0;
    endcase
  assign n7670 = n3006[1]; // extract
  assign n7671 = n5657[0]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7673 = 1'b0;
      13'b0100000000000: n7673 = 1'b0;
      13'b0010000000000: n7673 = n6878;
      13'b0001000000000: n7673 = 1'b0;
      13'b0000100000000: n7673 = 1'b0;
      13'b0000010000000: n7673 = 1'b0;
      13'b0000001000000: n7673 = 1'b0;
      13'b0000000100000: n7673 = 1'b0;
      13'b0000000010000: n7673 = 1'b0;
      13'b0000000001000: n7673 = 1'b0;
      13'b0000000000100: n7673 = n7671;
      13'b0000000000010: n7673 = 1'b0;
      13'b0000000000001: n7673 = n7670;
      default: n7673 = 1'b0;
    endcase
  assign n7674 = n3006[2]; // extract
  assign n7675 = n5657[1]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7677 = 1'b0;
      13'b0100000000000: n7677 = 1'b0;
      13'b0010000000000: n7677 = 1'b0;
      13'b0001000000000: n7677 = n6618;
      13'b0000100000000: n7677 = 1'b0;
      13'b0000010000000: n7677 = 1'b0;
      13'b0000001000000: n7677 = 1'b0;
      13'b0000000100000: n7677 = 1'b0;
      13'b0000000010000: n7677 = 1'b0;
      13'b0000000001000: n7677 = 1'b0;
      13'b0000000000100: n7677 = n7675;
      13'b0000000000010: n7677 = 1'b0;
      13'b0000000000001: n7677 = n7674;
      default: n7677 = 1'b0;
    endcase
  assign n7678 = n3006[3]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7680 = 1'b0;
      13'b0100000000000: n7680 = 1'b0;
      13'b0010000000000: n7680 = 1'b0;
      13'b0001000000000: n7680 = n6620;
      13'b0000100000000: n7680 = 1'b0;
      13'b0000010000000: n7680 = 1'b0;
      13'b0000001000000: n7680 = 1'b0;
      13'b0000000100000: n7680 = 1'b0;
      13'b0000000010000: n7680 = 1'b0;
      13'b0000000001000: n7680 = 1'b0;
      13'b0000000000100: n7680 = 1'b0;
      13'b0000000000010: n7680 = 1'b0;
      13'b0000000000001: n7680 = n7678;
      default: n7680 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7682 = 1'b0;
      13'b0100000000000: n7682 = n7274;
      13'b0010000000000: n7682 = 1'b0;
      13'b0001000000000: n7682 = 1'b0;
      13'b0000100000000: n7682 = 1'b0;
      13'b0000010000000: n7682 = 1'b0;
      13'b0000001000000: n7682 = 1'b0;
      13'b0000000100000: n7682 = 1'b0;
      13'b0000000010000: n7682 = 1'b0;
      13'b0000000001000: n7682 = 1'b0;
      13'b0000000000100: n7682 = 1'b0;
      13'b0000000000010: n7682 = 1'b0;
      13'b0000000000001: n7682 = 1'b0;
      default: n7682 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7684 = 1'b0;
      13'b0100000000000: n7684 = 1'b0;
      13'b0010000000000: n7684 = 1'b0;
      13'b0001000000000: n7684 = n6622;
      13'b0000100000000: n7684 = 1'b0;
      13'b0000010000000: n7684 = 1'b0;
      13'b0000001000000: n7684 = 1'b0;
      13'b0000000100000: n7684 = 1'b0;
      13'b0000000010000: n7684 = 1'b0;
      13'b0000000001000: n7684 = 1'b0;
      13'b0000000000100: n7684 = 1'b0;
      13'b0000000000010: n7684 = 1'b0;
      13'b0000000000001: n7684 = 1'b0;
      default: n7684 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7686 = 1'b0;
      13'b0100000000000: n7686 = 1'b0;
      13'b0010000000000: n7686 = 1'b0;
      13'b0001000000000: n7686 = 1'b0;
      13'b0000100000000: n7686 = 1'b0;
      13'b0000010000000: n7686 = 1'b0;
      13'b0000001000000: n7686 = 1'b0;
      13'b0000000100000: n7686 = 1'b0;
      13'b0000000010000: n7686 = 1'b0;
      13'b0000000001000: n7686 = 1'b0;
      13'b0000000000100: n7686 = n5658;
      13'b0000000000010: n7686 = 1'b0;
      13'b0000000000001: n7686 = 1'b0;
      default: n7686 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7688 = 1'b0;
      13'b0100000000000: n7688 = 1'b0;
      13'b0010000000000: n7688 = n6880;
      13'b0001000000000: n7688 = 1'b0;
      13'b0000100000000: n7688 = 1'b0;
      13'b0000010000000: n7688 = 1'b0;
      13'b0000001000000: n7688 = 1'b0;
      13'b0000000100000: n7688 = 1'b0;
      13'b0000000010000: n7688 = 1'b0;
      13'b0000000001000: n7688 = 1'b0;
      13'b0000000000100: n7688 = 1'b0;
      13'b0000000000010: n7688 = 1'b0;
      13'b0000000000001: n7688 = 1'b0;
      default: n7688 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7690 = 1'b0;
      13'b0100000000000: n7690 = 1'b0;
      13'b0010000000000: n7690 = 1'b0;
      13'b0001000000000: n7690 = 1'b0;
      13'b0000100000000: n7690 = 1'b0;
      13'b0000010000000: n7690 = 1'b0;
      13'b0000001000000: n7690 = n6295;
      13'b0000000100000: n7690 = 1'b0;
      13'b0000000010000: n7690 = 1'b0;
      13'b0000000001000: n7690 = 1'b0;
      13'b0000000000100: n7690 = n5660;
      13'b0000000000010: n7690 = 1'b0;
      13'b0000000000001: n7690 = 1'b0;
      default: n7690 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7692 = 1'b0;
      13'b0100000000000: n7692 = 1'b0;
      13'b0010000000000: n7692 = 1'b0;
      13'b0001000000000: n7692 = 1'b0;
      13'b0000100000000: n7692 = 1'b0;
      13'b0000010000000: n7692 = 1'b0;
      13'b0000001000000: n7692 = 1'b0;
      13'b0000000100000: n7692 = 1'b0;
      13'b0000000010000: n7692 = 1'b0;
      13'b0000000001000: n7692 = 1'b0;
      13'b0000000000100: n7692 = 1'b0;
      13'b0000000000010: n7692 = 1'b0;
      13'b0000000000001: n7692 = n3008;
      default: n7692 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7694 = 1'b0;
      13'b0100000000000: n7694 = 1'b0;
      13'b0010000000000: n7694 = 1'b0;
      13'b0001000000000: n7694 = 1'b0;
      13'b0000100000000: n7694 = 1'b0;
      13'b0000010000000: n7694 = 1'b0;
      13'b0000001000000: n7694 = 1'b0;
      13'b0000000100000: n7694 = 1'b0;
      13'b0000000010000: n7694 = 1'b0;
      13'b0000000001000: n7694 = 1'b0;
      13'b0000000000100: n7694 = n5662;
      13'b0000000000010: n7694 = 1'b0;
      13'b0000000000001: n7694 = 1'b0;
      default: n7694 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7696 = 1'b0;
      13'b0100000000000: n7696 = 1'b0;
      13'b0010000000000: n7696 = 1'b0;
      13'b0001000000000: n7696 = 1'b0;
      13'b0000100000000: n7696 = 1'b0;
      13'b0000010000000: n7696 = 1'b0;
      13'b0000001000000: n7696 = 1'b0;
      13'b0000000100000: n7696 = 1'b0;
      13'b0000000010000: n7696 = 1'b0;
      13'b0000000001000: n7696 = n5893;
      13'b0000000000100: n7696 = 1'b0;
      13'b0000000000010: n7696 = 1'b0;
      13'b0000000000001: n7696 = 1'b0;
      default: n7696 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7698 = 1'b0;
      13'b0100000000000: n7698 = 1'b0;
      13'b0010000000000: n7698 = n6882;
      13'b0001000000000: n7698 = 1'b0;
      13'b0000100000000: n7698 = 1'b0;
      13'b0000010000000: n7698 = 1'b0;
      13'b0000001000000: n7698 = 1'b0;
      13'b0000000100000: n7698 = 1'b0;
      13'b0000000010000: n7698 = 1'b0;
      13'b0000000001000: n7698 = 1'b0;
      13'b0000000000100: n7698 = 1'b0;
      13'b0000000000010: n7698 = 1'b0;
      13'b0000000000001: n7698 = 1'b0;
      default: n7698 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7700 = 1'b0;
      13'b0100000000000: n7700 = n7276;
      13'b0010000000000: n7700 = 1'b0;
      13'b0001000000000: n7700 = n6624;
      13'b0000100000000: n7700 = 1'b0;
      13'b0000010000000: n7700 = 1'b0;
      13'b0000001000000: n7700 = n6297;
      13'b0000000100000: n7700 = 1'b0;
      13'b0000000010000: n7700 = 1'b0;
      13'b0000000001000: n7700 = n5895;
      13'b0000000000100: n7700 = n5664;
      13'b0000000000010: n7700 = 1'b0;
      13'b0000000000001: n7700 = n3010;
      default: n7700 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7702 = 1'b0;
      13'b0100000000000: n7702 = 1'b0;
      13'b0010000000000: n7702 = 1'b0;
      13'b0001000000000: n7702 = 1'b0;
      13'b0000100000000: n7702 = 1'b0;
      13'b0000010000000: n7702 = 1'b0;
      13'b0000001000000: n7702 = 1'b0;
      13'b0000000100000: n7702 = 1'b0;
      13'b0000000010000: n7702 = 1'b0;
      13'b0000000001000: n7702 = 1'b0;
      13'b0000000000100: n7702 = n5666;
      13'b0000000000010: n7702 = 1'b0;
      13'b0000000000001: n7702 = 1'b0;
      default: n7702 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7704 = 1'b0;
      13'b0100000000000: n7704 = 1'b0;
      13'b0010000000000: n7704 = 1'b0;
      13'b0001000000000: n7704 = 1'b0;
      13'b0000100000000: n7704 = 1'b0;
      13'b0000010000000: n7704 = 1'b0;
      13'b0000001000000: n7704 = 1'b0;
      13'b0000000100000: n7704 = 1'b0;
      13'b0000000010000: n7704 = 1'b0;
      13'b0000000001000: n7704 = 1'b0;
      13'b0000000000100: n7704 = n5668;
      13'b0000000000010: n7704 = 1'b0;
      13'b0000000000001: n7704 = 1'b0;
      default: n7704 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7706 = 1'b0;
      13'b0100000000000: n7706 = 1'b0;
      13'b0010000000000: n7706 = 1'b0;
      13'b0001000000000: n7706 = 1'b0;
      13'b0000100000000: n7706 = 1'b0;
      13'b0000010000000: n7706 = 1'b0;
      13'b0000001000000: n7706 = 1'b0;
      13'b0000000100000: n7706 = 1'b0;
      13'b0000000010000: n7706 = 1'b0;
      13'b0000000001000: n7706 = 1'b0;
      13'b0000000000100: n7706 = n5670;
      13'b0000000000010: n7706 = 1'b0;
      13'b0000000000001: n7706 = 1'b0;
      default: n7706 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7708 = 2'b00;
      13'b0100000000000: n7708 = 2'b00;
      13'b0010000000000: n7708 = 2'b00;
      13'b0001000000000: n7708 = 2'b00;
      13'b0000100000000: n7708 = 2'b00;
      13'b0000010000000: n7708 = 2'b00;
      13'b0000001000000: n7708 = 2'b00;
      13'b0000000100000: n7708 = 2'b00;
      13'b0000000010000: n7708 = 2'b00;
      13'b0000000001000: n7708 = 2'b00;
      13'b0000000000100: n7708 = n5673;
      13'b0000000000010: n7708 = 2'b00;
      13'b0000000000001: n7708 = 2'b00;
      default: n7708 = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7710 = 1'b0;
      13'b0100000000000: n7710 = n7277;
      13'b0010000000000: n7710 = n6884;
      13'b0001000000000: n7710 = 1'b0;
      13'b0000100000000: n7710 = 1'b0;
      13'b0000010000000: n7710 = n6415;
      13'b0000001000000: n7710 = n6298;
      13'b0000000100000: n7710 = n5978;
      13'b0000000010000: n7710 = 1'b0;
      13'b0000000001000: n7710 = n5896;
      13'b0000000000100: n7710 = n5675;
      13'b0000000000010: n7710 = n3211;
      13'b0000000000001: n7710 = n3011;
      default: n7710 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7712 = 1'b0;
      13'b0100000000000: n7712 = 1'b0;
      13'b0010000000000: n7712 = n6886;
      13'b0001000000000: n7712 = 1'b0;
      13'b0000100000000: n7712 = 1'b0;
      13'b0000010000000: n7712 = 1'b0;
      13'b0000001000000: n7712 = 1'b0;
      13'b0000000100000: n7712 = 1'b0;
      13'b0000000010000: n7712 = 1'b0;
      13'b0000000001000: n7712 = 1'b0;
      13'b0000000000100: n7712 = 1'b0;
      13'b0000000000010: n7712 = 1'b0;
      13'b0000000000001: n7712 = 1'b0;
      default: n7712 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7714 = 2'b00;
      13'b0100000000000: n7714 = n7279;
      13'b0010000000000: n7714 = 2'b00;
      13'b0001000000000: n7714 = 2'b00;
      13'b0000100000000: n7714 = 2'b00;
      13'b0000010000000: n7714 = 2'b00;
      13'b0000001000000: n7714 = 2'b00;
      13'b0000000100000: n7714 = 2'b00;
      13'b0000000010000: n7714 = 2'b00;
      13'b0000000001000: n7714 = 2'b00;
      13'b0000000000100: n7714 = 2'b00;
      13'b0000000000010: n7714 = 2'b00;
      13'b0000000000001: n7714 = 2'b00;
      default: n7714 = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7716 = 2'b00;
      13'b0100000000000: n7716 = 2'b00;
      13'b0010000000000: n7716 = 2'b00;
      13'b0001000000000: n7716 = 2'b00;
      13'b0000100000000: n7716 = 2'b00;
      13'b0000010000000: n7716 = 2'b00;
      13'b0000001000000: n7716 = n6300;
      13'b0000000100000: n7716 = 2'b00;
      13'b0000000010000: n7716 = 2'b00;
      13'b0000000001000: n7716 = 2'b00;
      13'b0000000000100: n7716 = 2'b00;
      13'b0000000000010: n7716 = 2'b00;
      13'b0000000000001: n7716 = 2'b00;
      default: n7716 = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7718 = 1'b0;
      13'b0100000000000: n7718 = n7280;
      13'b0010000000000: n7718 = 1'b0;
      13'b0001000000000: n7718 = 1'b0;
      13'b0000100000000: n7718 = 1'b0;
      13'b0000010000000: n7718 = 1'b0;
      13'b0000001000000: n7718 = 1'b0;
      13'b0000000100000: n7718 = 1'b0;
      13'b0000000010000: n7718 = 1'b0;
      13'b0000000001000: n7718 = 1'b0;
      13'b0000000000100: n7718 = 1'b0;
      13'b0000000000010: n7718 = 1'b0;
      13'b0000000000001: n7718 = 1'b0;
      default: n7718 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7720 = 1'b0;
      13'b0100000000000: n7720 = 1'b0;
      13'b0010000000000: n7720 = 1'b0;
      13'b0001000000000: n7720 = 1'b0;
      13'b0000100000000: n7720 = 1'b0;
      13'b0000010000000: n7720 = 1'b0;
      13'b0000001000000: n7720 = 1'b0;
      13'b0000000100000: n7720 = 1'b0;
      13'b0000000010000: n7720 = 1'b0;
      13'b0000000001000: n7720 = 1'b0;
      13'b0000000000100: n7720 = n5676;
      13'b0000000000010: n7720 = 1'b0;
      13'b0000000000001: n7720 = 1'b0;
      default: n7720 = 1'b0;
    endcase
  assign n7740 = n7721[19:17]; // extract
  assign n7744 = n7721[27]; // extract
  assign n7746 = n7721[29]; // extract
  assign n7751 = n7721[66:35]; // extract
  assign n7753 = n7721[74:68]; // extract
  assign n7756 = n7721[80:79]; // extract
  assign n7757 = n7721[87:82]; // extract
  /* TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7425)
      13'b1000000000000: n7758 = n2057;
      13'b0100000000000: n7758 = n7281;
      13'b0010000000000: n7758 = n2057;
      13'b0001000000000: n7758 = n6625;
      13'b0000100000000: n7758 = n2057;
      13'b0000010000000: n7758 = n2057;
      13'b0000001000000: n7758 = n6301;
      13'b0000000100000: n7758 = n2057;
      13'b0000000010000: n7758 = n5955;
      13'b0000000001000: n7758 = n5897;
      13'b0000000000100: n7758 = n5677;
      13'b0000000000010: n7758 = n3178;
      13'b0000000000001: n7758 = n3012;
      default: n7758 = n2057;
    endcase
  /* TG68KdotC_Kernel.vhd:3186:36  */
  assign n7759 = set_exec[8]; // extract
  /* TG68KdotC_Kernel.vhd:3186:44  */
  assign n7760 = ~n7759;
  /* TG68KdotC_Kernel.vhd:3186:60  */
  assign n7761 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:3186:63  */
  assign n7762 = ~n7761;
  /* TG68KdotC_Kernel.vhd:3186:77  */
  assign n7763 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:3186:89  */
  assign n7765 = n7763 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3186:68  */
  assign n7766 = n7762 | n7765;
  /* TG68KdotC_Kernel.vhd:3186:49  */
  assign n7767 = n7766 & n7760;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7769 = n7791 ? 1'b1 : n7710;
  /* TG68KdotC_Kernel.vhd:3189:34  */
  assign n7770 = opcode[8]; // extract
  /* TG68KdotC_Kernel.vhd:3194:42  */
  assign n7772 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:3194:33  */
  assign n7774 = n7772 ? 1'b1 : n7453;
  /* TG68KdotC_Kernel.vhd:3197:33  */
  assign n7776 = setexecopc ? 1'b1 : n7471;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7778 = n7784 ? 1'b1 : n7440;
  /* TG68KdotC_Kernel.vhd:3189:25  */
  assign n7779 = n7770 ? n7453 : n7774;
  /* TG68KdotC_Kernel.vhd:3189:25  */
  assign n7781 = n7770 ? n7456 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3189:25  */
  assign n7782 = n7770 ? n7471 : n7776;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7783 = n7790 ? 1'b1 : n7700;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7784 = n7770 & build_logical;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7785 = build_logical ? n7779 : n7453;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7786 = build_logical ? n7781 : n7456;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7787 = build_logical ? n7782 : n7471;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7789 = build_logical ? 1'b1 : n7515;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7790 = n7770 & build_logical;
  /* TG68KdotC_Kernel.vhd:3184:17  */
  assign n7791 = n7767 & build_logical;
  /* TG68KdotC_Kernel.vhd:3209:34  */
  assign n7794 = opcode[3]; // extract
  /* TG68KdotC_Kernel.vhd:3211:50  */
  assign n7795 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:3211:62  */
  assign n7797 = n7795 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7799 = n7830 ? 1'b1 : n7572;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7803 = n7821 ? 2'b10 : n7430;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7805 = n7826 ? 1'b1 : n7465;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7806 = n7828 ? 1'b1 : n7544;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7807 = n7829 ? 1'b1 : n7564;
  /* TG68KdotC_Kernel.vhd:3210:33  */
  assign n7808 = n7797 & decodeopc;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7810 = n7834 ? 7'b0100001 : n7758;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7812 = decodeopc & n7794;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7813 = decodeopc & n7794;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7815 = n7794 ? n7787 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7816 = decodeopc & n7794;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7817 = decodeopc & n7794;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7818 = n7808 & n7794;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7819 = n7794 ? n7769 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3209:25  */
  assign n7820 = decodeopc & n7794;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7821 = n7812 & build_bcd;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7823 = build_bcd ? 1'b1 : n7778;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7825 = build_bcd ? 1'b1 : n7786;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7826 = n7813 & build_bcd;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7827 = build_bcd ? n7815 : n7787;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7828 = n7816 & build_bcd;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7829 = n7817 & build_bcd;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7830 = n7818 & build_bcd;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7831 = build_bcd ? 1'b1 : n7783;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7832 = build_bcd ? 1'b1 : n7702;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7833 = build_bcd ? n7819 : n7769;
  /* TG68KdotC_Kernel.vhd:3204:17  */
  assign n7834 = n7820 & build_bcd;
  /* TG68KdotC_Kernel.vhd:3231:33  */
  assign n7835 = ~trapd;
  /* TG68KdotC_Kernel.vhd:3229:17  */
  assign n7837 = n7838 ? 1'b1 : n7444;
  /* TG68KdotC_Kernel.vhd:3229:17  */
  assign n7838 = n7835 & set_z_error;
  /* TG68KdotC_Kernel.vhd:3229:17  */
  assign n7840 = set_z_error ? 1'b1 : n7509;
  /* TG68KdotC_Kernel.vhd:3242:25  */
  assign n7842 = clkena_lw ? trapmake : trapd;
  /* TG68KdotC_Kernel.vhd:3242:25  */
  assign n7843 = clkena_lw ? next_micro_state : micro_state;
  /* TG68KdotC_Kernel.vhd:3240:17  */
  assign n7844 = reset ? trapd : n7842;
  /* TG68KdotC_Kernel.vhd:3240:17  */
  assign n7846 = reset ? 7'b0000010 : n7843;
  /* TG68KdotC_Kernel.vhd:3249:33  */
  assign n7852 = micro_state == 7'b0000010;
  /* TG68KdotC_Kernel.vhd:3254:33  */
  assign n7855 = micro_state == 7'b0000011;
  /* TG68KdotC_Kernel.vhd:3259:33  */
  assign n7858 = micro_state == 7'b0000100;
  /* TG68KdotC_Kernel.vhd:3265:49  */
  assign n7859 = brief[8]; // extract
  /* TG68KdotC_Kernel.vhd:3265:52  */
  assign n7860 = ~n7859;
  /* TG68KdotC_Kernel.vhd:3265:57  */
  assign n7862 = n7860 | 1'b0;
  /* TG68KdotC_Kernel.vhd:3265:82  */
  assign n7863 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3265:85  */
  assign n7864 = ~n7863;
  /* TG68KdotC_Kernel.vhd:3265:90  */
  assign n7866 = 1'b1 & n7864;
  /* TG68KdotC_Kernel.vhd:3265:75  */
  assign n7867 = n7862 | n7866;
  /* TG68KdotC_Kernel.vhd:3272:57  */
  assign n7869 = brief[7]; // extract
  /* TG68KdotC_Kernel.vhd:3274:59  */
  assign n7870 = exec[22]; // extract
  /* TG68KdotC_Kernel.vhd:3274:49  */
  assign n7872 = n7870 ? 1'b1 : n2041;
  /* TG68KdotC_Kernel.vhd:3272:49  */
  assign n7874 = n7869 ? 1'b1 : n2034;
  /* TG68KdotC_Kernel.vhd:3272:49  */
  assign n7875 = n7869 ? n2041 : n7872;
  /* TG68KdotC_Kernel.vhd:3277:57  */
  assign n7876 = brief[5]; // extract
  /* TG68KdotC_Kernel.vhd:3277:60  */
  assign n7877 = ~n7876;
  /* TG68KdotC_Kernel.vhd:3280:65  */
  assign n7878 = brief[4]; // extract
  /* TG68KdotC_Kernel.vhd:3280:57  */
  assign n7880 = n7878 ? 1'b1 : n7601;
  /* TG68KdotC_Kernel.vhd:3277:49  */
  assign n7882 = n7877 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3277:49  */
  assign n7883 = n7877 ? n7601 : n7880;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7885 = n7867 ? 2'b01 : n7882;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7888 = n7867 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7891 = n7867 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7892 = n7867 ? n2034 : n7874;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7893 = n7867 ? n2041 : n7875;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7894 = n7867 ? 1'b1 : n7643;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7895 = n7867 ? n7601 : n7883;
  /* TG68KdotC_Kernel.vhd:3265:41  */
  assign n7898 = n7867 ? 7'b0000110 : 7'b0001011;
  /* TG68KdotC_Kernel.vhd:3264:33  */
  assign n7900 = micro_state == 7'b0000101;
  /* TG68KdotC_Kernel.vhd:3287:33  */
  assign n7903 = micro_state == 7'b0000110;
  /* TG68KdotC_Kernel.vhd:3295:49  */
  assign n7904 = brief[5]; // extract
  /* TG68KdotC_Kernel.vhd:3295:41  */
  assign n7907 = n7904 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3298:49  */
  assign n7908 = brief[6]; // extract
  /* TG68KdotC_Kernel.vhd:3298:52  */
  assign n7909 = ~n7908;
  /* TG68KdotC_Kernel.vhd:3298:66  */
  assign n7910 = brief[2]; // extract
  /* TG68KdotC_Kernel.vhd:3298:69  */
  assign n7911 = ~n7910;
  /* TG68KdotC_Kernel.vhd:3298:57  */
  assign n7912 = n7911 & n7909;
  /* TG68KdotC_Kernel.vhd:3301:57  */
  assign n7914 = brief[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:3301:69  */
  assign n7916 = n7914 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3301:49  */
  assign n7919 = n7916 ? 7'b0000110 : 7'b0001100;
  /* TG68KdotC_Kernel.vhd:3307:57  */
  assign n7920 = brief[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:3307:69  */
  assign n7922 = n7920 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3307:49  */
  assign n7926 = n7922 ? n7803 : 2'b10;
  /* TG68KdotC_Kernel.vhd:3307:49  */
  assign n7929 = n7922 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3307:49  */
  assign n7931 = n7922 ? 1'b1 : n7431;
  /* TG68KdotC_Kernel.vhd:3307:49  */
  assign n7932 = n7922 ? 1'b1 : n2047;
  /* TG68KdotC_Kernel.vhd:3307:49  */
  assign n7933 = n7922 ? n7601 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3307:49  */
  assign n7935 = n7922 ? n7810 : 7'b0001101;
  /* TG68KdotC_Kernel.vhd:3298:41  */
  assign n7937 = n7912 ? 2'b01 : n7926;
  /* TG68KdotC_Kernel.vhd:3298:41  */
  assign n7939 = n7912 ? 1'b0 : n7929;
  /* TG68KdotC_Kernel.vhd:3298:41  */
  assign n7940 = n7912 ? n7431 : n7931;
  /* TG68KdotC_Kernel.vhd:3298:41  */
  assign n7941 = n7912 ? n2047 : n7932;
  /* TG68KdotC_Kernel.vhd:3298:41  */
  assign n7942 = n7912 ? 1'b1 : n7643;
  /* TG68KdotC_Kernel.vhd:3298:41  */
  assign n7943 = n7912 ? n7601 : n7933;
  /* TG68KdotC_Kernel.vhd:3298:41  */
  assign n7944 = n7912 ? n7919 : n7935;
  /* TG68KdotC_Kernel.vhd:3294:33  */
  assign n7946 = micro_state == 7'b0001011;
  /* TG68KdotC_Kernel.vhd:3318:33  */
  assign n7949 = micro_state == 7'b0001100;
  /* TG68KdotC_Kernel.vhd:3328:49  */
  assign n7951 = brief[1]; // extract
  /* TG68KdotC_Kernel.vhd:3328:52  */
  assign n7952 = ~n7951;
  /* TG68KdotC_Kernel.vhd:3331:57  */
  assign n7953 = brief[0]; // extract
  /* TG68KdotC_Kernel.vhd:3331:49  */
  assign n7955 = n7953 ? 1'b1 : n7601;
  /* TG68KdotC_Kernel.vhd:3328:41  */
  assign n7957 = n7952 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3328:41  */
  assign n7958 = n7952 ? n7601 : n7955;
  /* TG68KdotC_Kernel.vhd:3325:33  */
  assign n7960 = micro_state == 7'b0001101;
  /* TG68KdotC_Kernel.vhd:3338:49  */
  assign n7961 = brief[1]; // extract
  /* TG68KdotC_Kernel.vhd:3338:41  */
  assign n7964 = n7961 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3341:49  */
  assign n7965 = brief[6]; // extract
  /* TG68KdotC_Kernel.vhd:3341:52  */
  assign n7966 = ~n7965;
  /* TG68KdotC_Kernel.vhd:3341:66  */
  assign n7967 = brief[2]; // extract
  /* TG68KdotC_Kernel.vhd:3341:57  */
  assign n7968 = n7967 & n7966;
  /* TG68KdotC_Kernel.vhd:3341:41  */
  assign n7972 = n7968 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3341:41  */
  assign n7974 = n7968 ? n7431 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3341:41  */
  assign n7975 = n7968 ? n2047 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3341:41  */
  assign n7976 = n7968 ? 1'b1 : n7643;
  /* TG68KdotC_Kernel.vhd:3341:41  */
  assign n7978 = n7968 ? 7'b0000110 : n7810;
  /* TG68KdotC_Kernel.vhd:3337:33  */
  assign n7980 = micro_state == 7'b0001110;
  /* TG68KdotC_Kernel.vhd:3351:33  */
  assign n7982 = micro_state == 7'b0000111;
  /* TG68KdotC_Kernel.vhd:3357:49  */
  assign n7983 = brief[8]; // extract
  /* TG68KdotC_Kernel.vhd:3357:52  */
  assign n7984 = ~n7983;
  /* TG68KdotC_Kernel.vhd:3357:57  */
  assign n7986 = n7984 | 1'b0;
  /* TG68KdotC_Kernel.vhd:3357:82  */
  assign n7987 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3357:85  */
  assign n7988 = ~n7987;
  /* TG68KdotC_Kernel.vhd:3357:90  */
  assign n7990 = 1'b1 & n7988;
  /* TG68KdotC_Kernel.vhd:3357:75  */
  assign n7991 = n7986 | n7990;
  /* TG68KdotC_Kernel.vhd:3364:57  */
  assign n7993 = brief[7]; // extract
  /* TG68KdotC_Kernel.vhd:3364:49  */
  assign n7995 = n7993 ? 1'b1 : n2034;
  /* TG68KdotC_Kernel.vhd:3369:57  */
  assign n7996 = brief[5]; // extract
  /* TG68KdotC_Kernel.vhd:3369:60  */
  assign n7997 = ~n7996;
  /* TG68KdotC_Kernel.vhd:3372:65  */
  assign n7998 = brief[4]; // extract
  /* TG68KdotC_Kernel.vhd:3372:57  */
  assign n8000 = n7998 ? 1'b1 : n7601;
  /* TG68KdotC_Kernel.vhd:3369:49  */
  assign n8002 = n7997 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3369:49  */
  assign n8003 = n7997 ? n7601 : n8000;
  /* TG68KdotC_Kernel.vhd:3357:41  */
  assign n8005 = n7991 ? 2'b01 : n8002;
  /* TG68KdotC_Kernel.vhd:3357:41  */
  assign n8008 = n7991 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3357:41  */
  assign n8011 = n7991 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3357:41  */
  assign n8012 = n7991 ? n2034 : n7995;
  /* TG68KdotC_Kernel.vhd:3357:41  */
  assign n8013 = n7991 ? 1'b1 : n7643;
  /* TG68KdotC_Kernel.vhd:3357:41  */
  assign n8014 = n7991 ? n7601 : n8003;
  /* TG68KdotC_Kernel.vhd:3357:41  */
  assign n8017 = n7991 ? 7'b0010100 : 7'b0001111;
  /* TG68KdotC_Kernel.vhd:3356:33  */
  assign n8019 = micro_state == 7'b0010011;
  /* TG68KdotC_Kernel.vhd:3379:33  */
  assign n8022 = micro_state == 7'b0010100;
  /* TG68KdotC_Kernel.vhd:3388:49  */
  assign n8023 = brief[5]; // extract
  /* TG68KdotC_Kernel.vhd:3388:41  */
  assign n8026 = n8023 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3391:49  */
  assign n8027 = brief[6]; // extract
  /* TG68KdotC_Kernel.vhd:3391:52  */
  assign n8028 = ~n8027;
  /* TG68KdotC_Kernel.vhd:3391:66  */
  assign n8029 = brief[2]; // extract
  /* TG68KdotC_Kernel.vhd:3391:69  */
  assign n8030 = ~n8029;
  /* TG68KdotC_Kernel.vhd:3391:57  */
  assign n8031 = n8030 & n8028;
  /* TG68KdotC_Kernel.vhd:3394:57  */
  assign n8033 = brief[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:3394:69  */
  assign n8035 = n8033 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3394:49  */
  assign n8038 = n8035 ? 7'b0010100 : 7'b0010000;
  /* TG68KdotC_Kernel.vhd:3400:57  */
  assign n8039 = brief[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:3400:69  */
  assign n8041 = n8039 == 2'b00;
  /* TG68KdotC_Kernel.vhd:3400:49  */
  assign n8046 = n8041 ? 2'b11 : 2'b10;
  assign n8047 = n7595[1]; // extract
  /* TG68KdotC_Kernel.vhd:3400:49  */
  assign n8048 = n8041 ? n8047 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3400:49  */
  assign n8049 = n8041 ? n7601 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3400:49  */
  assign n8052 = n8041 ? 7'b0000001 : 7'b0010001;
  /* TG68KdotC_Kernel.vhd:3391:41  */
  assign n8054 = n8031 ? 2'b01 : n8046;
  assign n8055 = n7595[1]; // extract
  /* TG68KdotC_Kernel.vhd:3391:41  */
  assign n8056 = n8031 ? n8055 : n8048;
  /* TG68KdotC_Kernel.vhd:3391:41  */
  assign n8057 = n8031 ? 1'b1 : n7643;
  /* TG68KdotC_Kernel.vhd:3391:41  */
  assign n8058 = n8031 ? n7601 : n8049;
  /* TG68KdotC_Kernel.vhd:3391:41  */
  assign n8059 = n8031 ? n8038 : n8052;
  /* TG68KdotC_Kernel.vhd:3387:33  */
  assign n8061 = micro_state == 7'b0001111;
  /* TG68KdotC_Kernel.vhd:3411:33  */
  assign n8065 = micro_state == 7'b0010000;
  /* TG68KdotC_Kernel.vhd:3422:49  */
  assign n8068 = brief[1]; // extract
  /* TG68KdotC_Kernel.vhd:3422:52  */
  assign n8069 = ~n8068;
  /* TG68KdotC_Kernel.vhd:3425:57  */
  assign n8070 = brief[0]; // extract
  /* TG68KdotC_Kernel.vhd:3425:49  */
  assign n8072 = n8070 ? 1'b1 : n7601;
  /* TG68KdotC_Kernel.vhd:3422:41  */
  assign n8074 = n8069 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3422:41  */
  assign n8075 = n8069 ? n7601 : n8072;
  /* TG68KdotC_Kernel.vhd:3418:33  */
  assign n8077 = micro_state == 7'b0010001;
  /* TG68KdotC_Kernel.vhd:3433:49  */
  assign n8079 = brief[1]; // extract
  /* TG68KdotC_Kernel.vhd:3433:41  */
  assign n8082 = n8079 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3436:49  */
  assign n8083 = brief[6]; // extract
  /* TG68KdotC_Kernel.vhd:3436:52  */
  assign n8084 = ~n8083;
  /* TG68KdotC_Kernel.vhd:3436:66  */
  assign n8085 = brief[2]; // extract
  /* TG68KdotC_Kernel.vhd:3436:57  */
  assign n8086 = n8085 & n8084;
  /* TG68KdotC_Kernel.vhd:3436:41  */
  assign n8090 = n8086 ? 2'b01 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3436:41  */
  assign n8091 = n8086 ? 1'b1 : n7643;
  /* TG68KdotC_Kernel.vhd:3436:41  */
  assign n8094 = n8086 ? 7'b0010100 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3431:33  */
  assign n8096 = micro_state == 7'b0010010;
  /* TG68KdotC_Kernel.vhd:3447:41  */
  assign n8098 = exe_condition ? 1'b1 : n7426;
  /* TG68KdotC_Kernel.vhd:3447:41  */
  assign n8101 = exe_condition ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3447:41  */
  assign n8103 = exe_condition ? 7'b0000001 : n7810;
  /* TG68KdotC_Kernel.vhd:3446:33  */
  assign n8105 = micro_state == 7'b0010101;
  /* TG68KdotC_Kernel.vhd:3453:33  */
  assign n8107 = micro_state == 7'b0010110;
  /* TG68KdotC_Kernel.vhd:3458:54  */
  assign n8108 = ~long_start;
  /* TG68KdotC_Kernel.vhd:3458:41  */
  assign n8111 = n8108 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3457:33  */
  assign n8114 = micro_state == 7'b0010111;
  /* TG68KdotC_Kernel.vhd:3467:33  */
  assign n8116 = micro_state == 7'b0011000;
  /* TG68KdotC_Kernel.vhd:3471:57  */
  assign n8117 = ~exe_condition;
  /* TG68KdotC_Kernel.vhd:3473:57  */
  assign n8118 = c_out[1]; // extract
  /* TG68KdotC_Kernel.vhd:3471:41  */
  assign n8120 = n8126 ? 1'b1 : n7426;
  /* TG68KdotC_Kernel.vhd:3473:49  */
  assign n8123 = n8118 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3471:41  */
  assign n8125 = n8132 ? 7'b0000001 : n7810;
  /* TG68KdotC_Kernel.vhd:3471:41  */
  assign n8126 = n8118 & n8117;
  /* TG68KdotC_Kernel.vhd:3471:41  */
  assign n8129 = n8117 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3471:41  */
  assign n8131 = n8117 ? n8123 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3471:41  */
  assign n8132 = n8118 & n8117;
  /* TG68KdotC_Kernel.vhd:3470:33  */
  assign n8134 = micro_state == 7'b0011001;
  /* TG68KdotC_Kernel.vhd:3480:33  */
  assign n8140 = micro_state == 7'b1000001;
  /* TG68KdotC_Kernel.vhd:3489:50  */
  assign n8141 = sndopc[15]; // extract
  /* TG68KdotC_Kernel.vhd:3492:58  */
  assign n8142 = opcode[10:9]; // extract
  /* TG68KdotC_Kernel.vhd:3492:71  */
  assign n8144 = n8142 == 2'b00;
  assign n8146 = n1788[88]; // extract
  /* TG68KdotC_Kernel.vhd:3489:41  */
  assign n8147 = n8154 ? 1'b1 : n8146;
  /* TG68KdotC_Kernel.vhd:3489:41  */
  assign n8149 = n8141 ? 2'b10 : n7429;
  /* TG68KdotC_Kernel.vhd:3489:41  */
  assign n8152 = n8141 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3489:41  */
  assign n8154 = n8144 & n8141;
  /* TG68KdotC_Kernel.vhd:3487:33  */
  assign n8159 = micro_state == 7'b1000010;
  /* TG68KdotC_Kernel.vhd:3504:50  */
  assign n8161 = sndopc[15]; // extract
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8163 = n8161 ? 2'b10 : n7429;
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8166 = n8161 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3511:61  */
  assign n8170 = exec[88]; // extract
  /* TG68KdotC_Kernel.vhd:3512:50  */
  assign n8171 = sndopc[11]; // extract
  /* TG68KdotC_Kernel.vhd:3512:41  */
  assign n8173 = n8171 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3512:41  */
  assign n8175 = n8171 ? 7'b1000100 : n7810;
  /* TG68KdotC_Kernel.vhd:3501:33  */
  assign n8177 = micro_state == 7'b1000011;
  /* TG68KdotC_Kernel.vhd:3516:33  */
  assign n8179 = micro_state == 7'b1000100;
  /* TG68KdotC_Kernel.vhd:3520:49  */
  assign n8180 = flags[0]; // extract
  /* TG68KdotC_Kernel.vhd:3520:41  */
  assign n8182 = n8180 ? 1'b1 : n7840;
  /* TG68KdotC_Kernel.vhd:3519:33  */
  assign n8184 = micro_state == 7'b1000101;
  /* TG68KdotC_Kernel.vhd:3525:33  */
  assign n8186 = micro_state == 7'b0110111;
  /* TG68KdotC_Kernel.vhd:3530:49  */
  assign n8187 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8194 = n8187 ? 2'b11 : n7803;
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8197 = n8187 ? 1'b0 : 1'b1;
  assign n8198 = n1788[27]; // extract
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8199 = n8187 ? n8198 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8200 = n8187 ? n7539 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8201 = n8187 ? 1'b1 : n7548;
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8202 = n8187 ? 1'b1 : n1804;
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8203 = n8187 ? n7612 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3530:41  */
  assign n8205 = n8187 ? 7'b0000001 : n7810;
  /* TG68KdotC_Kernel.vhd:3528:33  */
  assign n8207 = micro_state == 7'b0111000;
  /* TG68KdotC_Kernel.vhd:3544:63  */
  assign n8208 = sndopc[15]; // extract
  /* TG68KdotC_Kernel.vhd:3542:33  */
  assign n8211 = micro_state == 7'b0111001;
  /* TG68KdotC_Kernel.vhd:3547:33  */
  assign n8217 = micro_state == 7'b0111010;
  /* TG68KdotC_Kernel.vhd:3555:33  */
  assign n8220 = micro_state == 7'b0111011;
  /* TG68KdotC_Kernel.vhd:3560:49  */
  assign n8221 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:3560:41  */
  assign n8223 = n8221 ? 1'b1 : n7614;
  /* TG68KdotC_Kernel.vhd:3559:33  */
  assign n8229 = micro_state == 7'b0111100;
  /* TG68KdotC_Kernel.vhd:3570:33  */
  assign n8232 = micro_state == 7'b0111101;
  /* TG68KdotC_Kernel.vhd:3575:49  */
  assign n8233 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:3579:71  */
  assign n8235 = sndopc[15]; // extract
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8243 = n8233 ? 2'b11 : n7803;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8246 = n8233 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8248 = n8233 ? n8235 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8251 = n8233 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8253 = n8233 ? 1'b1 : n7468;
  assign n8254 = n1788[27]; // extract
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8255 = n8233 ? n8254 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8256 = n8233 ? n7539 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8257 = n8233 ? 1'b1 : n7548;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8258 = n8233 ? 1'b1 : n2047;
  assign n8259 = n7595[1]; // extract
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8260 = n8233 ? n8259 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8261 = n8233 ? n7608 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8262 = n8233 ? n7612 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8265 = n8233 ? 7'b0111111 : 7'b1000000;
  /* TG68KdotC_Kernel.vhd:3574:33  */
  assign n8267 = micro_state == 7'b0111110;
  /* TG68KdotC_Kernel.vhd:3592:33  */
  assign n8271 = micro_state == 7'b0111111;
  /* TG68KdotC_Kernel.vhd:3599:33  */
  assign n8275 = micro_state == 7'b1000000;
  /* TG68KdotC_Kernel.vhd:3605:58  */
  assign n8276 = last_data_read[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:3605:71  */
  assign n8278 = n8276 != 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3607:58  */
  assign n8279 = opcode[5:3]; // extract
  /* TG68KdotC_Kernel.vhd:3607:70  */
  assign n8281 = n8279 == 3'b100;
  /* TG68KdotC_Kernel.vhd:3609:63  */
  assign n8283 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3605:41  */
  assign n8285 = n8290 ? 1'b1 : n7539;
  /* TG68KdotC_Kernel.vhd:3607:49  */
  assign n8286 = n8283 & n8281;
  /* TG68KdotC_Kernel.vhd:3605:41  */
  assign n8287 = n8291 ? 1'b1 : n7585;
  /* TG68KdotC_Kernel.vhd:3605:41  */
  assign n8289 = n8278 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3605:41  */
  assign n8290 = n8286 & n8278;
  /* TG68KdotC_Kernel.vhd:3605:41  */
  assign n8291 = n8281 & n8278;
  /* TG68KdotC_Kernel.vhd:3605:41  */
  assign n8293 = n8278 ? 7'b0011011 : n7810;
  /* TG68KdotC_Kernel.vhd:3604:33  */
  assign n8295 = micro_state == 7'b0011010;
  /* TG68KdotC_Kernel.vhd:3616:53  */
  assign n8296 = ~movem_run;
  /* TG68KdotC_Kernel.vhd:3622:58  */
  assign n8299 = opcode[10]; // extract
  /* TG68KdotC_Kernel.vhd:3622:62  */
  assign n8300 = ~n8299;
  /* TG68KdotC_Kernel.vhd:3622:49  */
  assign n8304 = n8300 ? 2'b11 : 2'b10;
  /* TG68KdotC_Kernel.vhd:3622:49  */
  assign n8305 = n8300 ? 1'b1 : n7548;
  /* TG68KdotC_Kernel.vhd:3616:41  */
  assign n8307 = n8296 ? 2'b01 : n8304;
  /* TG68KdotC_Kernel.vhd:3616:41  */
  assign n8308 = n8296 ? n7548 : n8305;
  /* TG68KdotC_Kernel.vhd:3616:41  */
  assign n8309 = n8296 ? n7585 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3616:41  */
  assign n8310 = n8296 ? n7597 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3616:41  */
  assign n8312 = n8296 ? n7810 : 7'b0011011;
  /* TG68KdotC_Kernel.vhd:3615:33  */
  assign n8314 = micro_state == 7'b0011011;
  /* TG68KdotC_Kernel.vhd:3631:50  */
  assign n8315 = opcode[5:4]; // extract
  /* TG68KdotC_Kernel.vhd:3631:62  */
  assign n8317 = n8315 != 2'b00;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8319 = n8317 ? 1'b1 : n7431;
  /* TG68KdotC_Kernel.vhd:3630:33  */
  assign n8321 = micro_state == 7'b0011101;
  /* TG68KdotC_Kernel.vhd:3636:50  */
  assign n8322 = opcode[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:3636:62  */
  assign n8324 = n8322 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3636:41  */
  assign n8326 = n8324 ? 1'b1 : n7799;
  /* TG68KdotC_Kernel.vhd:3635:33  */
  assign n8331 = micro_state == 7'b0011110;
  /* TG68KdotC_Kernel.vhd:3646:50  */
  assign n8332 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3646:63  */
  assign n8334 = n8332 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3646:41  */
  assign n8336 = n8334 ? 1'b1 : n7799;
  /* TG68KdotC_Kernel.vhd:3651:50  */
  assign n8338 = opcode[7:6]; // extract
  /* TG68KdotC_Kernel.vhd:3651:63  */
  assign n8340 = n8338 == 2'b01;
  /* TG68KdotC_Kernel.vhd:3651:41  */
  assign n8343 = n8340 ? 2'b00 : 2'b01;
  /* TG68KdotC_Kernel.vhd:3645:33  */
  assign n8346 = micro_state == 7'b0011111;
  /* TG68KdotC_Kernel.vhd:3661:33  */
  assign n8348 = micro_state == 7'b0100000;
  /* TG68KdotC_Kernel.vhd:3665:50  */
  assign n8349 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3665:63  */
  assign n8351 = n8349 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3665:41  */
  assign n8353 = n8351 ? 1'b1 : n7799;
  /* TG68KdotC_Kernel.vhd:3664:33  */
  assign n8356 = micro_state == 7'b0100001;
  /* TG68KdotC_Kernel.vhd:3675:50  */
  assign n8357 = opcode[11:9]; // extract
  /* TG68KdotC_Kernel.vhd:3675:63  */
  assign n8359 = n8357 == 3'b111;
  /* TG68KdotC_Kernel.vhd:3675:41  */
  assign n8361 = n8359 ? 1'b1 : n7799;
  /* TG68KdotC_Kernel.vhd:3674:33  */
  assign n8364 = micro_state == 7'b0100010;
  /* TG68KdotC_Kernel.vhd:3684:33  */
  assign n8368 = micro_state == 7'b0100011;
  /* TG68KdotC_Kernel.vhd:3690:33  */
  assign n8371 = micro_state == 7'b0100100;
  /* TG68KdotC_Kernel.vhd:3694:33  */
  assign n8374 = micro_state == 7'b0100101;
  /* TG68KdotC_Kernel.vhd:3699:33  */
  assign n8377 = micro_state == 7'b0100110;
  /* TG68KdotC_Kernel.vhd:3703:33  */
  assign n8380 = micro_state == 7'b0110010;
  /* TG68KdotC_Kernel.vhd:3720:71  */
  assign n8383 = trap_interrupt | trap_trace;
  /* TG68KdotC_Kernel.vhd:3720:89  */
  assign n8384 = n8383 | trap_berr;
  /* TG68KdotC_Kernel.vhd:3720:49  */
  assign n8386 = n8384 ? 1'b1 : n7837;
  /* TG68KdotC_Kernel.vhd:3714:41  */
  assign n8389 = use_vbr_stackframe ? 2'b01 : 2'b10;
  /* TG68KdotC_Kernel.vhd:3714:41  */
  assign n8390 = use_vbr_stackframe ? n7837 : n8386;
  /* TG68KdotC_Kernel.vhd:3714:41  */
  assign n8391 = use_vbr_stackframe ? 1'b1 : n1837;
  /* TG68KdotC_Kernel.vhd:3714:41  */
  assign n8394 = use_vbr_stackframe ? 7'b0110100 : 7'b0110101;
  /* TG68KdotC_Kernel.vhd:3710:33  */
  assign n8396 = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:3728:63  */
  assign n8397 = trap_interrupt | trap_trace;
  /* TG68KdotC_Kernel.vhd:3728:41  */
  assign n8399 = n8397 ? 1'b1 : n7837;
  /* TG68KdotC_Kernel.vhd:3727:33  */
  assign n8402 = micro_state == 7'b0110100;
  /* TG68KdotC_Kernel.vhd:3742:41  */
  assign n8406 = trap_berr ? 7'b1000110 : 7'b0110110;
  /* TG68KdotC_Kernel.vhd:3736:33  */
  assign n8408 = micro_state == 7'b0110101;
  /* TG68KdotC_Kernel.vhd:3747:33  */
  assign n8412 = micro_state == 7'b0110110;
  /* TG68KdotC_Kernel.vhd:3754:33  */
  assign n8415 = micro_state == 7'b1000110;
  /* TG68KdotC_Kernel.vhd:3761:33  */
  assign n8418 = micro_state == 7'b1000111;
  /* TG68KdotC_Kernel.vhd:3768:33  */
  assign n8421 = micro_state == 7'b1001000;
  /* TG68KdotC_Kernel.vhd:3789:62  */
  assign n8424 = ~use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:3789:76  */
  assign n8425 = opcode[2]; // extract
  /* TG68KdotC_Kernel.vhd:3789:67  */
  assign n8426 = n8424 | n8425;
  /* TG68KdotC_Kernel.vhd:3789:41  */
  assign n8429 = n8426 ? 1'b1 : n7626;
  assign n8430 = n7590[1]; // extract
  /* TG68KdotC_Kernel.vhd:3789:41  */
  assign n8431 = n8426 ? 1'b1 : n8430;
  /* TG68KdotC_Kernel.vhd:3783:33  */
  assign n8433 = micro_state == 7'b0101011;
  /* TG68KdotC_Kernel.vhd:3797:77  */
  assign n8435 = opcode[2]; // extract
  /* TG68KdotC_Kernel.vhd:3797:80  */
  assign n8436 = ~n8435;
  /* TG68KdotC_Kernel.vhd:3797:67  */
  assign n8437 = n8436 & use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:3797:41  */
  assign n8440 = n8437 ? 2'b10 : n7803;
  /* TG68KdotC_Kernel.vhd:3797:41  */
  assign n8442 = n8437 ? 1'b1 : n7442;
  /* TG68KdotC_Kernel.vhd:3797:41  */
  assign n8443 = n8437 ? 1'b1 : n7560;
  /* TG68KdotC_Kernel.vhd:3797:41  */
  assign n8446 = n8437 ? 7'b0101101 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3794:33  */
  assign n8448 = micro_state == 7'b0101100;
  /* TG68KdotC_Kernel.vhd:3810:33  */
  assign n8450 = micro_state == 7'b0101101;
  /* TG68KdotC_Kernel.vhd:3817:56  */
  assign n8451 = last_data_in[15:12]; // extract
  /* TG68KdotC_Kernel.vhd:3817:70  */
  assign n8453 = n8451 == 4'b0010;
  /* TG68KdotC_Kernel.vhd:3817:41  */
  assign n8457 = n8453 ? 2'b10 : 2'b01;
  /* TG68KdotC_Kernel.vhd:3817:41  */
  assign n8459 = n8453 ? 2'b10 : n7803;
  /* TG68KdotC_Kernel.vhd:3817:41  */
  assign n8461 = n8453 ? 1'b1 : n7442;
  /* TG68KdotC_Kernel.vhd:3817:41  */
  assign n8462 = n8453 ? 1'b1 : n7560;
  /* TG68KdotC_Kernel.vhd:3817:41  */
  assign n8465 = n8453 ? 7'b0101111 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3815:33  */
  assign n8467 = micro_state == 7'b0101110;
  /* TG68KdotC_Kernel.vhd:3828:33  */
  assign n8469 = micro_state == 7'b0101111;
  /* TG68KdotC_Kernel.vhd:3832:33  */
  assign n8471 = micro_state == 7'b0110000;
  /* TG68KdotC_Kernel.vhd:3834:33  */
  assign n8474 = micro_state == 7'b0110001;
  /* TG68KdotC_Kernel.vhd:3841:50  */
  assign n8476 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3841:63  */
  assign n8478 = n8476 == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:3841:79  */
  assign n8479 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3841:92  */
  assign n8481 = n8479 == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:3841:71  */
  assign n8482 = n8478 | n8481;
  /* TG68KdotC_Kernel.vhd:3841:108  */
  assign n8483 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3841:121  */
  assign n8485 = n8483 == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:3841:100  */
  assign n8486 = n8482 | n8485;
  /* TG68KdotC_Kernel.vhd:3841:137  */
  assign n8487 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3841:150  */
  assign n8489 = n8487 == 12'b100000000001;
  /* TG68KdotC_Kernel.vhd:3841:129  */
  assign n8490 = n8486 | n8489;
  /* TG68KdotC_Kernel.vhd:3842:48  */
  assign n8491 = CPU[1]; // extract
  /* TG68KdotC_Kernel.vhd:3842:66  */
  assign n8492 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3842:79  */
  assign n8494 = n8492 == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:3842:95  */
  assign n8495 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3842:108  */
  assign n8497 = n8495 == 12'b100000000010;
  /* TG68KdotC_Kernel.vhd:3842:87  */
  assign n8498 = n8494 | n8497;
  /* TG68KdotC_Kernel.vhd:3842:124  */
  assign n8499 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3842:137  */
  assign n8501 = n8499 == 12'b100000000011;
  /* TG68KdotC_Kernel.vhd:3842:116  */
  assign n8502 = n8498 | n8501;
  /* TG68KdotC_Kernel.vhd:3842:153  */
  assign n8503 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:3842:166  */
  assign n8505 = n8503 == 12'b100000000100;
  /* TG68KdotC_Kernel.vhd:3842:145  */
  assign n8506 = n8502 | n8505;
  /* TG68KdotC_Kernel.vhd:3842:56  */
  assign n8507 = n8506 & n8491;
  /* TG68KdotC_Kernel.vhd:3841:159  */
  assign n8508 = n8490 | n8507;
  /* TG68KdotC_Kernel.vhd:3843:58  */
  assign n8509 = opcode[0]; // extract
  /* TG68KdotC_Kernel.vhd:3843:61  */
  assign n8510 = ~n8509;
  /* TG68KdotC_Kernel.vhd:3841:41  */
  assign n8512 = n8517 ? 1'b1 : n7539;
  /* TG68KdotC_Kernel.vhd:3841:41  */
  assign n8514 = n8508 ? n7487 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3841:41  */
  assign n8516 = n8508 ? n7840 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3841:41  */
  assign n8517 = n8510 & n8508;
  /* TG68KdotC_Kernel.vhd:3838:33  */
  assign n8519 = micro_state == 7'b1001001;
  /* TG68KdotC_Kernel.vhd:3859:50  */
  assign n8523 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:3859:41  */
  assign n8525 = n8523 ? 1'b1 : n7543;
  /* TG68KdotC_Kernel.vhd:3862:50  */
  assign n8526 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:3862:53  */
  assign n8527 = ~n8526;
  /* TG68KdotC_Kernel.vhd:3862:41  */
  assign n8530 = n8527 ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3854:33  */
  assign n8532 = micro_state == 7'b1001010;
  /* TG68KdotC_Kernel.vhd:3869:50  */
  assign n8533 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:3869:41  */
  assign n8536 = n8533 ? 1'b1 : n7546;
  /* TG68KdotC_Kernel.vhd:3869:41  */
  assign n8537 = n8533 ? 1'b1 : n7585;
  /* TG68KdotC_Kernel.vhd:3873:50  */
  assign n8538 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:3873:53  */
  assign n8539 = ~n8538;
  /* TG68KdotC_Kernel.vhd:3873:41  */
  assign n8542 = n8539 ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3868:33  */
  assign n8544 = micro_state == 7'b1001011;
  /* TG68KdotC_Kernel.vhd:3880:50  */
  assign n8545 = opcode[6]; // extract
  /* TG68KdotC_Kernel.vhd:3884:58  */
  assign n8549 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:3884:61  */
  assign n8550 = ~n8549;
  /* TG68KdotC_Kernel.vhd:3884:49  */
  assign n8553 = n8550 ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3880:41  */
  assign n8555 = n8545 ? n7428 : 2'b01;
  /* TG68KdotC_Kernel.vhd:3880:41  */
  assign n8556 = n8545 ? n8553 : n7803;
  /* TG68KdotC_Kernel.vhd:3880:41  */
  assign n8557 = n8545 ? 1'b1 : n7546;
  /* TG68KdotC_Kernel.vhd:3880:41  */
  assign n8558 = n8545 ? 1'b1 : n7585;
  /* TG68KdotC_Kernel.vhd:3880:41  */
  assign n8559 = n8545 ? 1'b1 : n7642;
  /* TG68KdotC_Kernel.vhd:3880:41  */
  assign n8561 = n8545 ? 7'b1001101 : n7810;
  /* TG68KdotC_Kernel.vhd:3879:33  */
  assign n8563 = micro_state == 7'b1001100;
  /* TG68KdotC_Kernel.vhd:3894:50  */
  assign n8564 = opcode[7]; // extract
  /* TG68KdotC_Kernel.vhd:3894:53  */
  assign n8565 = ~n8564;
  /* TG68KdotC_Kernel.vhd:3894:41  */
  assign n8568 = n8565 ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3893:33  */
  assign n8570 = micro_state == 7'b1001101;
  /* TG68KdotC_Kernel.vhd:3900:33  */
  assign n8572 = micro_state == 7'b1001110;
  /* TG68KdotC_Kernel.vhd:3904:50  */
  assign n8573 = opcode[15]; // extract
  /* TG68KdotC_Kernel.vhd:3904:59  */
  assign n8575 = n8573 | 1'b0;
  /* TG68KdotC_Kernel.vhd:3904:41  */
  assign n8578 = n8575 ? 6'b001110 : 6'b011110;
  /* TG68KdotC_Kernel.vhd:3903:33  */
  assign n8580 = micro_state == 7'b1010001;
  /* TG68KdotC_Kernel.vhd:3913:51  */
  assign n8583 = rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:3913:41  */
  assign n8586 = n8583 ? 7'b1010011 : 7'b1010010;
  /* TG68KdotC_Kernel.vhd:3911:33  */
  assign n8588 = micro_state == 7'b1010010;
  /* TG68KdotC_Kernel.vhd:3920:50  */
  assign n8589 = opcode[15]; // extract
  /* TG68KdotC_Kernel.vhd:3920:54  */
  assign n8590 = ~n8589;
  /* TG68KdotC_Kernel.vhd:3920:41  */
  assign n8592 = n8590 ? 1'b1 : n7608;
  /* TG68KdotC_Kernel.vhd:3925:50  */
  assign n8594 = opcode[15]; // extract
  /* TG68KdotC_Kernel.vhd:3925:54  */
  assign n8595 = ~n8594;
  /* TG68KdotC_Kernel.vhd:3925:59  */
  assign n8597 = 1'b1 & n8595;
  /* TG68KdotC_Kernel.vhd:3928:58  */
  assign n8599 = sndopc[10]; // extract
  /* TG68KdotC_Kernel.vhd:3925:41  */
  assign n8601 = n8605 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3925:41  */
  assign n8603 = n8611 ? 7'b1010100 : n7810;
  /* TG68KdotC_Kernel.vhd:3925:41  */
  assign n8605 = n8599 & n8597;
  /* TG68KdotC_Kernel.vhd:3925:41  */
  assign n8607 = n8597 ? 1'b1 : n7468;
  /* TG68KdotC_Kernel.vhd:3925:41  */
  assign n8608 = n8597 ? 1'b1 : n7539;
  assign n8609 = n7595[4]; // extract
  /* TG68KdotC_Kernel.vhd:3925:41  */
  assign n8610 = n8597 ? 1'b1 : n8609;
  /* TG68KdotC_Kernel.vhd:3925:41  */
  assign n8611 = n8599 & n8597;
  /* TG68KdotC_Kernel.vhd:3919:33  */
  assign n8613 = micro_state == 7'b1010011;
  /* TG68KdotC_Kernel.vhd:3935:33  */
  assign n8618 = micro_state == 7'b1010100;
  /* TG68KdotC_Kernel.vhd:3941:33  */
  assign n8620 = micro_state == 7'b1010101;
  /* TG68KdotC_Kernel.vhd:3945:51  */
  assign n8621 = op2out[31:16]; // extract
  /* TG68KdotC_Kernel.vhd:3945:65  */
  assign n8623 = n8621 == 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3945:83  */
  assign n8624 = opcode[15]; // extract
  /* TG68KdotC_Kernel.vhd:3945:74  */
  assign n8625 = n8623 | n8624;
  /* TG68KdotC_Kernel.vhd:3945:92  */
  assign n8627 = n8625 | 1'b0;
  /* TG68KdotC_Kernel.vhd:3945:117  */
  assign n8628 = op2out[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:3945:130  */
  assign n8630 = n8628 == 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3945:107  */
  assign n8631 = n8630 & n8627;
  /* TG68KdotC_Kernel.vhd:3945:41  */
  assign n8634 = n8631 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3945:41  */
  assign n8636 = n8631 ? n7810 : 7'b1010111;
  /* TG68KdotC_Kernel.vhd:3944:33  */
  assign n8639 = micro_state == 7'b1010110;
  /* TG68KdotC_Kernel.vhd:3953:50  */
  assign n8640 = opcode[15]; // extract
  /* TG68KdotC_Kernel.vhd:3953:59  */
  assign n8642 = n8640 | 1'b0;
  /* TG68KdotC_Kernel.vhd:3953:41  */
  assign n8645 = n8642 ? 6'b001101 : 6'b011101;
  /* TG68KdotC_Kernel.vhd:3952:33  */
  assign n8647 = micro_state == 7'b1010111;
  /* TG68KdotC_Kernel.vhd:3962:51  */
  assign n8650 = rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8653 = n8650 ? 7'b1011001 : 7'b1011000;
  /* TG68KdotC_Kernel.vhd:3960:33  */
  assign n8655 = micro_state == 7'b1011000;
  /* TG68KdotC_Kernel.vhd:3968:51  */
  assign n8656 = ~z_error;
  /* TG68KdotC_Kernel.vhd:3968:70  */
  assign n8657 = ~set_v_flag;
  /* TG68KdotC_Kernel.vhd:3968:56  */
  assign n8658 = n8657 & n8656;
  /* TG68KdotC_Kernel.vhd:3968:41  */
  assign n8660 = n8658 ? 1'b1 : n7539;
  /* TG68KdotC_Kernel.vhd:3971:50  */
  assign n8661 = opcode[15]; // extract
  /* TG68KdotC_Kernel.vhd:3971:54  */
  assign n8662 = ~n8661;
  /* TG68KdotC_Kernel.vhd:3971:59  */
  assign n8664 = 1'b1 & n8662;
  /* TG68KdotC_Kernel.vhd:3971:41  */
  assign n8667 = n8664 ? 2'b01 : n7803;
  /* TG68KdotC_Kernel.vhd:3971:41  */
  assign n8670 = n8664 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3971:41  */
  assign n8671 = n8664 ? 1'b1 : n7641;
  /* TG68KdotC_Kernel.vhd:3971:41  */
  assign n8673 = n8664 ? 7'b1011010 : n7810;
  /* TG68KdotC_Kernel.vhd:3967:33  */
  assign n8676 = micro_state == 7'b1011001;
  /* TG68KdotC_Kernel.vhd:3980:48  */
  assign n8677 = exec[34]; // extract
  /* TG68KdotC_Kernel.vhd:3980:41  */
  assign n8680 = n8677 ? 1'b1 : n7539;
  /* TG68KdotC_Kernel.vhd:3980:41  */
  assign n8681 = n8677 ? n7570 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3979:33  */
  assign n8684 = micro_state == 7'b1011010;
  /* TG68KdotC_Kernel.vhd:3989:50  */
  assign n8685 = op2out[5:0]; // extract
  /* TG68KdotC_Kernel.vhd:3989:62  */
  assign n8687 = n8685 != 6'b000000;
  /* TG68KdotC_Kernel.vhd:3990:70  */
  assign n8688 = op2out[5:0]; // extract
  assign n8690 = {n7479, n7476};
  /* TG68KdotC_Kernel.vhd:3989:41  */
  assign n8691 = n8687 ? n8688 : n8690;
  assign n8692 = n7721[23]; // extract
  /* TG68KdotC_Kernel.vhd:3989:41  */
  assign n8693 = n8687 ? n8692 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3988:33  */
  assign n8695 = micro_state == 7'b1001111;
  /* TG68KdotC_Kernel.vhd:3995:33  */
  assign n8697 = micro_state == 7'b1010000;
  assign n8698 = {n8697, n8695, n8684, n8676, n8655, n8647, n8639, n8620, n8618, n8613, n8588, n8580, n8572, n8570, n8563, n8544, n8532, n8519, n8474, n8471, n8469, n8467, n8450, n8448, n8433, n8421, n8418, n8415, n8412, n8408, n8402, n8396, n8380, n8377, n8374, n8371, n8368, n8364, n8356, n8348, n8346, n8331, n8321, n8314, n8295, n8275, n8271, n8267, n8232, n8229, n8220, n8217, n8211, n8207, n8186, n8184, n8179, n8177, n8159, n8140, n8134, n8116, n8114, n8107, n8105, n8096, n8077, n8065, n8061, n8022, n8019, n7982, n7980, n7960, n7949, n7946, n7903, n7900, n7858, n7855, n7852};
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8701 = 1'b1;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8701 = n8120;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8701 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8701 = n8098;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8701 = n7426;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8701 = n7426;
      default: n8701 = n7426;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8714 = n8555;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8714 = n8457;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8714 = 2'b01;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8714 = 2'b01;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8714 = 2'b01;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8714 = 2'b01;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8714 = n8389;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8714 = 2'b10;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8714 = n8343;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8714 = n7428;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8714 = n7428;
      default: n8714 = n7428;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8715 = n8163;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8715 = n8149;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8715 = n7429;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8715 = n7429;
      default: n8715 = n7429;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = n8667;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = 2'b01;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = 2'b01;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = 2'b01;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = 2'b01;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8753 = n8601;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8753 = 2'b01;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8753 = 2'b01;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8753 = n8568;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8753 = n8556;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8753 = n8542;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8753 = n8530;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8753 = n8459;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8753 = n8440;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8753 = 2'b10;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8753 = n8307;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8753 = n8289;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8753 = n8243;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8753 = n8194;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8753 = n8173;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8753 = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8753 = n8090;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8753 = n8074;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8753 = 2'b10;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8753 = n8054;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8753 = n8005;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8753 = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8753 = n7972;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8753 = n7957;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8753 = 2'b10;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8753 = n7937;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8753 = n7885;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8753 = n7803;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8753 = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8753 = n7803;
      default: n8753 = n7803;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8756 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8756 = n7939;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8756 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8756 = 1'b0;
      default: n8756 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8759 = n8129;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8759 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8759 = 1'b0;
      default: n8759 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8764 = n8319;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8764 = n7974;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8764 = n7940;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8764 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8764 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8764 = n7431;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8764 = 1'b1;
      default: n8764 = n7431;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8766 = n8008;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8766 = n7888;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8766 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8766 = 1'b0;
      default: n8766 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8776 = n8082;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8776 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8776 = n8026;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8776 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8776 = n8011;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8776 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8776 = n7964;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8776 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8776 = n7907;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8776 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8776 = n7891;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8776 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8776 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8776 = 1'b0;
      default: n8776 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8780 = n8131;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8780 = n8111;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8780 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8780 = n8101;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8780 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8780 = 1'b0;
      default: n8780 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8794 = n8461;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8794 = n8442;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8794 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8794 = n7442;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8794 = n7442;
      default: n8794 = n7442;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8796 = n8399;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8796 = n8390;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8796 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8796 = n7837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8796 = n7837;
      default: n8796 = n7837;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b1;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8799 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8799 = 1'b0;
      default: n8799 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8802 = 1'b1;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8802 = n7785;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8802 = n7785;
      default: n8802 = n7785;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8805 = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8805 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8805 = 1'b0;
      default: n8805 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8809 = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8809 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8809 = 1'b0;
      default: n8809 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8813 = n8246;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8813 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8813 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8813 = 1'b0;
      default: n8813 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8816 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8816 = n7462;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8816 = n7462;
      default: n8816 = n7462;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8821 = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8821 = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8821 = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8821 = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8821 = n7805;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8821 = n7805;
      default: n8821 = n7805;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8823 = n8248;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8823 = n8208;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8823 = n8166;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8823 = n8152;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8823 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8823 = 1'b0;
      default: n8823 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8828 = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8828 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8828 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8828 = 1'b0;
      default: n8828 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8831 = n8251;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8831 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8831 = 1'b0;
      default: n8831 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = 1'b1;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n8607;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8837 = n8253;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8837 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8837 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8837 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8837 = n7468;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8837 = n7468;
      default: n8837 = n7468;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = n8670;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8841 = 1'b1;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8841 = n8197;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8841 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8841 = 1'b0;
      default: n8841 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8846 = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8846 = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8846 = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8846 = n7827;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8846 = n7827;
      default: n8846 = n7827;
    endcase
  assign n8847 = {n7479, n7476};
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8691;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8645;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8578;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8848 = n8847;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8848 = n8847;
      default: n8848 = n8847;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8852 = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8852 = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8852 = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8852 = n7484;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8852 = n7484;
      default: n8852 = n7484;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8855 = 1'b1;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8855 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8855 = 1'b0;
      default: n8855 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8862 = 1'b1;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8862 = 1'b1;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8862 = 1'b1;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8862 = 1'b1;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8862 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8862 = 1'b0;
      default: n8862 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8864 = n8514;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8864 = n7487;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8864 = n7487;
      default: n8864 = n7487;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8865 = n8516;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8865 = n8182;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8865 = n7840;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8865 = n7840;
      default: n8865 = n7840;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8868 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8868 = n8012;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8868 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8868 = n7892;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8868 = n2034;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8868 = n2034;
      default: n8868 = n2034;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = n8634;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8870 = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8870 = 1'b0;
      default: n8870 = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8872 = 1'b1;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8872 = n7527;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8872 = n7527;
      default: n8872 = n7527;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8873 = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8873 = 1'b1;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8873 = n7531;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8873 = n7531;
      default: n8873 = n7531;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = 1'b1;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = 1'b1;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8874 = n7618;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8874 = n7618;
      default: n8874 = n7618;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8875 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8875 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8875 = n7893;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8875 = n2041;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8875 = n2041;
      default: n8875 = n2041;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = 1'b1;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8876 = n7533;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8876 = n7533;
      default: n8876 = n7533;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8877 = n8391;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8877 = n1837;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8877 = n1837;
      default: n8877 = n1837;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8878 = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8878 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8878 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8878 = n7535;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8878 = n7535;
      default: n8878 = n7535;
    endcase
  assign n8879 = n1788[27]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8880 = 1'b1;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8880 = 1'b1;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8880 = n8255;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8880 = n8199;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8880 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8880 = n8879;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8880 = n8879;
      default: n8880 = n8879;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n8680;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n8660;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8881 = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n8608;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8881 = n8512;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8881 = 1'b1;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8881 = 1'b1;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8881 = n8285;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8881 = 1'b1;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8881 = n8256;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8881 = n8200;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8881 = n7539;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8881 = n7539;
      default: n8881 = n7539;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8882 = 1'b1;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8882 = n8429;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8882 = n7626;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8882 = n7626;
      default: n8882 = n7626;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8883 = n8525;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8883 = n7543;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8883 = n7543;
      default: n8883 = n7543;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8884 = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8884 = n7806;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8884 = n7806;
      default: n8884 = n7806;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8885 = n8557;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8885 = n8536;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8885 = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8885 = n7546;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8885 = n7546;
      default: n8885 = n7546;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8886 = n8308;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8886 = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8886 = n8257;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8886 = n8201;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8886 = n7548;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8886 = n7548;
      default: n8886 = n7548;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8887 = n7630;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8887 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8887 = 1'b1;
      default: n8887 = n7630;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8888 = n8462;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8888 = n8443;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8888 = 1'b1;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8888 = 1'b1;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8888 = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8888 = n7560;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8888 = n7560;
      default: n8888 = n7560;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8889 = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8889 = n7807;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8889 = n7807;
      default: n8889 = n7807;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n8681;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8890 = n7570;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8890 = n7570;
      default: n8890 = n7570;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8891 = n8361;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8891 = n8353;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8891 = n8336;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8891 = n8326;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8891 = n7799;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8891 = n7799;
      default: n8891 = n7799;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8892 = n8558;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8892 = n8537;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8892 = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8892 = n8309;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8892 = n8287;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8892 = n7585;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8892 = n7585;
      default: n8892 = n7585;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8893 = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8893 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8893 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8893 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8893 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8893 = n7588;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8893 = n7588;
      default: n8893 = n7588;
    endcase
  assign n8894 = n7590[0]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8895 = 1'b1;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8895 = 1'b1;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8895 = n8894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8895 = n8894;
      default: n8895 = n8894;
    endcase
  assign n8896 = n7590[1]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8897 = n8431;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8897 = 1'b1;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8897 = n8896;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8897 = n8896;
      default: n8897 = n8896;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8898 = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8898 = n8258;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8898 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8898 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8898 = n7975;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8898 = n7941;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8898 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8898 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8898 = n2047;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8898 = 1'b1;
      default: n8898 = n2047;
    endcase
  assign n8899 = n7595[1]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8900 = n8260;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8900 = 1'b1;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8900 = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8900 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8900 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8900 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8900 = n8056;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8900 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8900 = n8899;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8900 = n8899;
      default: n8900 = n8899;
    endcase
  assign n8901 = n7595[4]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8610;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8902 = n8901;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8902 = n8901;
      default: n8902 = n8901;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n8671;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8903 = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8903 = n7641;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8903 = n7641;
      default: n8903 = n7641;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8904 = n8310;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8904 = n7597;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8904 = n7597;
      default: n8904 = n7597;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8905 = 1'b1;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8905 = n8091;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8905 = n8057;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8905 = n8013;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8905 = n7976;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8905 = n7942;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8905 = n7894;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8905 = n7643;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8905 = n7643;
      default: n8905 = n7643;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8906 = n8559;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8906 = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8906 = n7642;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8906 = n7642;
      default: n8906 = n7642;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8907 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8907 = n8075;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8907 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8907 = n8058;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8907 = n8014;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8907 = n7958;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8907 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8907 = n7943;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8907 = n7895;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8907 = n7601;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8907 = n7601;
      default: n8907 = n7601;
    endcase
  assign n8908 = n1788[79]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8909 = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8909 = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8909 = n8908;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8909 = n8908;
      default: n8909 = n8908;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n8592;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8910 = n8261;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8910 = n7608;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8910 = n7608;
      default: n8910 = n7608;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8911 = n8202;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8911 = n1804;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8911 = n1804;
      default: n8911 = n1804;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8912 = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8912 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8912 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8912 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8912 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8912 = n7610;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8912 = n7610;
      default: n8912 = n7610;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8913 = 1'b1;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8913 = n8262;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8913 = n8203;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8913 = n7612;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8913 = n7612;
      default: n8913 = n7612;
    endcase
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8914 = n8223;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8914 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8914 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8914 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8914 = n7614;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8914 = n7614;
      default: n8914 = n7614;
    endcase
  assign n8915 = n1788[87]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8916 = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8916 = n8915;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8916 = n8915;
      default: n8916 = n8915;
    endcase
  assign n8917 = n1788[88]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8918 = n8170;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8918 = n8147;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8918 = n8917;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8918 = n8917;
      default: n8918 = n8917;
    endcase
  assign n8919 = n1788[28]; // extract
  assign n8921 = n7590[3:2]; // extract
  assign n8923 = n7595[0]; // extract
  assign n8924 = n7595[3:2]; // extract
  assign n8925 = n1788[78:75]; // extract
  assign n8927 = n7721[23]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8693;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8928 = n8927;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8928 = n8927;
      default: n8928 = n8927;
    endcase
  assign n8929 = n7721[25:24]; // extract
  assign n8930 = n7721[22:21]; // extract
  /* TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8698)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n8673;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n8653;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b1011000;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n8636;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b1010110;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n8603;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8971 = n8586;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b1010010;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b1001110;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8971 = n8561;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b1001100;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b1001011;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b0110001;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8971 = 7'b0000001;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8971 = n8465;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8971 = 7'b0101110;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8971 = n8446;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8971 = 7'b0101100;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8971 = 7'b0110110;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8971 = 7'b1001000;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8971 = 7'b1000111;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8971 = 7'b0011000;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8971 = n8406;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8971 = 7'b0110101;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8971 = n8394;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8971 = 7'b0110011;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8971 = 7'b0100110;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8971 = 7'b0100100;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8971 = 7'b0100000;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8971 = 7'b0011111;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8971 = n8312;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8971 = n8293;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8971 = 7'b0011000;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8971 = n8265;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8971 = 7'b0111110;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8971 = 7'b0111101;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8971 = 7'b0111100;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8971 = 7'b0111011;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8971 = 7'b0111010;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8971 = n8205;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8971 = 7'b0111000;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8971 = n7810;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8971 = 7'b1000101;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8971 = n8175;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8971 = 7'b1000011;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8971 = 7'b1000010;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8971 = n8125;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8971 = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8971 = 7'b0011000;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8971 = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8971 = n8103;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8971 = n8094;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8971 = 7'b0010010;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8971 = 7'b0010001;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8971 = n8059;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8971 = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8971 = n8017;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8971 = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8971 = n7978;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8971 = 7'b0001110;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8971 = 7'b0001101;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8971 = n7944;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8971 = n7810;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8971 = n7898;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8971 = n7810;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8971 = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8971 = n7810;
      default: n8971 = n7810;
    endcase
  /* TG68KdotC_Kernel.vhd:4012:41  */
  assign n8977 = exec[33]; // extract
  /* TG68KdotC_Kernel.vhd:4012:33  */
  assign n8978 = n8977 & clkena_lw;
  /* TG68KdotC_Kernel.vhd:4013:27  */
  assign n8979 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:4014:47  */
  assign n8980 = reg_qa[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:4014:19  */
  assign n8982 = n8979 == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:4015:47  */
  assign n8983 = reg_qa[2:0]; // extract
  /* TG68KdotC_Kernel.vhd:4015:19  */
  assign n8985 = n8979 == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:4016:48  */
  assign n8986 = reg_qa[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:4016:19  */
  assign n8988 = n8979 == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:4017:19  */
  assign n8990 = n8979 == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:4018:19  */
  assign n8992 = n8979 == 12'b100000000001;
  /* TG68KdotC_Kernel.vhd:4019:19  */
  assign n8994 = n8979 == 12'b100000000010;
  /* TG68KdotC_Kernel.vhd:4020:19  */
  assign n8996 = n8979 == 12'b100000000011;
  /* TG68KdotC_Kernel.vhd:4021:19  */
  assign n8998 = n8979 == 12'b100000000100;
  assign n8999 = {n8998, n8996, n8994, n8992, n8990, n8988, n8985, n8982};
  /* TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n8999)
      8'b10000000: n9000 = vbr;
      8'b01000000: n9000 = vbr;
      8'b00100000: n9000 = vbr;
      8'b00010000: n9000 = reg_qa;
      8'b00001000: n9000 = vbr;
      8'b00000100: n9000 = vbr;
      8'b00000010: n9000 = vbr;
      8'b00000001: n9000 = vbr;
      default: n9000 = vbr;
    endcase
  /* TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n8999)
      8'b10000000: n9001 = cacr;
      8'b01000000: n9001 = cacr;
      8'b00100000: n9001 = cacr;
      8'b00010000: n9001 = cacr;
      8'b00001000: n9001 = cacr;
      8'b00000100: n9001 = n8986;
      8'b00000010: n9001 = cacr;
      8'b00000001: n9001 = cacr;
      default: n9001 = cacr;
    endcase
  /* TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n8999)
      8'b10000000: n9002 = dfc;
      8'b01000000: n9002 = dfc;
      8'b00100000: n9002 = dfc;
      8'b00010000: n9002 = dfc;
      8'b00001000: n9002 = dfc;
      8'b00000100: n9002 = dfc;
      8'b00000010: n9002 = n8983;
      8'b00000001: n9002 = dfc;
      default: n9002 = dfc;
    endcase
  /* TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n8999)
      8'b10000000: n9003 = sfc;
      8'b01000000: n9003 = sfc;
      8'b00100000: n9003 = sfc;
      8'b00010000: n9003 = sfc;
      8'b00001000: n9003 = sfc;
      8'b00000100: n9003 = sfc;
      8'b00000010: n9003 = sfc;
      8'b00000001: n9003 = n8980;
      default: n9003 = sfc;
    endcase
  /* TG68KdotC_Kernel.vhd:4012:11  */
  assign n9004 = n8978 ? n9000 : vbr;
  /* TG68KdotC_Kernel.vhd:4012:11  */
  assign n9005 = n8978 ? n9001 : cacr;
  /* TG68KdotC_Kernel.vhd:4012:11  */
  assign n9006 = n8978 ? n9002 : dfc;
  /* TG68KdotC_Kernel.vhd:4012:11  */
  assign n9007 = n8978 ? n9003 : sfc;
  /* TG68KdotC_Kernel.vhd:4009:11  */
  assign n9009 = reset ? 32'b00000000000000000000000000000000 : n9004;
  /* TG68KdotC_Kernel.vhd:4009:11  */
  assign n9011 = reset ? 4'b0000 : n9005;
  /* TG68KdotC_Kernel.vhd:4009:11  */
  assign n9012 = reset ? dfc : n9006;
  /* TG68KdotC_Kernel.vhd:4009:11  */
  assign n9013 = reset ? sfc : n9007;
  /* TG68KdotC_Kernel.vhd:4028:19  */
  assign n9018 = brief[11:0]; // extract
  /* TG68KdotC_Kernel.vhd:4029:78  */
  assign n9020 = {29'b00000000000000000000000000000, sfc};
  /* TG68KdotC_Kernel.vhd:4029:17  */
  assign n9022 = n9018 == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:4030:78  */
  assign n9024 = {29'b00000000000000000000000000000, dfc};
  /* TG68KdotC_Kernel.vhd:4030:17  */
  assign n9026 = n9018 == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:4031:79  */
  assign n9028 = cacr & 4'b0011;
  /* TG68KdotC_Kernel.vhd:4031:71  */
  assign n9030 = {28'b0000000000000000000000000000, n9028};
  /* TG68KdotC_Kernel.vhd:4031:11  */
  assign n9032 = n9018 == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:4033:11  */
  assign n9034 = n9018 == 12'b100000000001;
  assign n9035 = {n9034, n9032, n9026, n9022};
  /* TG68KdotC_Kernel.vhd:4028:9  */
  always @*
    case (n9035)
      4'b1000: n9037 = vbr;
      4'b0100: n9037 = n9030;
      4'b0010: n9037 = n9024;
      4'b0001: n9037 = n9020;
      default: n9037 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68KdotC_Kernel.vhd:4047:32  */
  assign n9042 = exe_opcode[11:8]; // extract
  /* TG68KdotC_Kernel.vhd:4048:25  */
  assign n9044 = n9042 == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4049:25  */
  assign n9046 = n9042 == 4'b0001;
  /* TG68KdotC_Kernel.vhd:4050:65  */
  assign n9047 = flags[0]; // extract
  /* TG68KdotC_Kernel.vhd:4050:56  */
  assign n9048 = ~n9047;
  /* TG68KdotC_Kernel.vhd:4050:82  */
  assign n9049 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:4050:73  */
  assign n9050 = ~n9049;
  /* TG68KdotC_Kernel.vhd:4050:69  */
  assign n9051 = n9048 & n9050;
  /* TG68KdotC_Kernel.vhd:4050:25  */
  assign n9053 = n9042 == 4'b0010;
  /* TG68KdotC_Kernel.vhd:4051:60  */
  assign n9054 = flags[0]; // extract
  /* TG68KdotC_Kernel.vhd:4051:72  */
  assign n9055 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:4051:64  */
  assign n9056 = n9054 | n9055;
  /* TG68KdotC_Kernel.vhd:4051:25  */
  assign n9058 = n9042 == 4'b0011;
  /* TG68KdotC_Kernel.vhd:4052:64  */
  assign n9059 = flags[0]; // extract
  /* TG68KdotC_Kernel.vhd:4052:55  */
  assign n9060 = ~n9059;
  /* TG68KdotC_Kernel.vhd:4052:25  */
  assign n9062 = n9042 == 4'b0100;
  /* TG68KdotC_Kernel.vhd:4053:60  */
  assign n9063 = flags[0]; // extract
  /* TG68KdotC_Kernel.vhd:4053:25  */
  assign n9065 = n9042 == 4'b0101;
  /* TG68KdotC_Kernel.vhd:4054:64  */
  assign n9066 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:4054:55  */
  assign n9067 = ~n9066;
  /* TG68KdotC_Kernel.vhd:4054:25  */
  assign n9069 = n9042 == 4'b0110;
  /* TG68KdotC_Kernel.vhd:4055:60  */
  assign n9070 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:4055:25  */
  assign n9072 = n9042 == 4'b0111;
  /* TG68KdotC_Kernel.vhd:4056:64  */
  assign n9073 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4056:55  */
  assign n9074 = ~n9073;
  /* TG68KdotC_Kernel.vhd:4056:25  */
  assign n9076 = n9042 == 4'b1000;
  /* TG68KdotC_Kernel.vhd:4057:60  */
  assign n9077 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4057:25  */
  assign n9079 = n9042 == 4'b1001;
  /* TG68KdotC_Kernel.vhd:4058:64  */
  assign n9080 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4058:55  */
  assign n9081 = ~n9080;
  /* TG68KdotC_Kernel.vhd:4058:25  */
  assign n9083 = n9042 == 4'b1010;
  /* TG68KdotC_Kernel.vhd:4059:60  */
  assign n9084 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4059:25  */
  assign n9086 = n9042 == 4'b1011;
  /* TG68KdotC_Kernel.vhd:4060:61  */
  assign n9087 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4060:74  */
  assign n9088 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4060:65  */
  assign n9089 = n9087 & n9088;
  /* TG68KdotC_Kernel.vhd:4060:92  */
  assign n9090 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4060:83  */
  assign n9091 = ~n9090;
  /* TG68KdotC_Kernel.vhd:4060:109  */
  assign n9092 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4060:100  */
  assign n9093 = ~n9092;
  /* TG68KdotC_Kernel.vhd:4060:96  */
  assign n9094 = n9091 & n9093;
  /* TG68KdotC_Kernel.vhd:4060:79  */
  assign n9095 = n9089 | n9094;
  /* TG68KdotC_Kernel.vhd:4060:25  */
  assign n9097 = n9042 == 4'b1100;
  /* TG68KdotC_Kernel.vhd:4061:61  */
  assign n9098 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4061:78  */
  assign n9099 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4061:69  */
  assign n9100 = ~n9099;
  /* TG68KdotC_Kernel.vhd:4061:65  */
  assign n9101 = n9098 & n9100;
  /* TG68KdotC_Kernel.vhd:4061:96  */
  assign n9102 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4061:87  */
  assign n9103 = ~n9102;
  /* TG68KdotC_Kernel.vhd:4061:109  */
  assign n9104 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4061:100  */
  assign n9105 = n9103 & n9104;
  /* TG68KdotC_Kernel.vhd:4061:83  */
  assign n9106 = n9101 | n9105;
  /* TG68KdotC_Kernel.vhd:4061:25  */
  assign n9108 = n9042 == 4'b1101;
  /* TG68KdotC_Kernel.vhd:4062:61  */
  assign n9109 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4062:74  */
  assign n9110 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4062:65  */
  assign n9111 = n9109 & n9110;
  /* TG68KdotC_Kernel.vhd:4062:91  */
  assign n9112 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:4062:82  */
  assign n9113 = ~n9112;
  /* TG68KdotC_Kernel.vhd:4062:78  */
  assign n9114 = n9111 & n9113;
  /* TG68KdotC_Kernel.vhd:4062:109  */
  assign n9115 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4062:100  */
  assign n9116 = ~n9115;
  /* TG68KdotC_Kernel.vhd:4062:126  */
  assign n9117 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4062:117  */
  assign n9118 = ~n9117;
  /* TG68KdotC_Kernel.vhd:4062:113  */
  assign n9119 = n9116 & n9118;
  /* TG68KdotC_Kernel.vhd:4062:143  */
  assign n9120 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:4062:134  */
  assign n9121 = ~n9120;
  /* TG68KdotC_Kernel.vhd:4062:130  */
  assign n9122 = n9119 & n9121;
  /* TG68KdotC_Kernel.vhd:4062:96  */
  assign n9123 = n9114 | n9122;
  /* TG68KdotC_Kernel.vhd:4062:25  */
  assign n9125 = n9042 == 4'b1110;
  /* TG68KdotC_Kernel.vhd:4063:61  */
  assign n9126 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4063:78  */
  assign n9127 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4063:69  */
  assign n9128 = ~n9127;
  /* TG68KdotC_Kernel.vhd:4063:65  */
  assign n9129 = n9126 & n9128;
  /* TG68KdotC_Kernel.vhd:4063:96  */
  assign n9130 = flags[3]; // extract
  /* TG68KdotC_Kernel.vhd:4063:87  */
  assign n9131 = ~n9130;
  /* TG68KdotC_Kernel.vhd:4063:109  */
  assign n9132 = flags[1]; // extract
  /* TG68KdotC_Kernel.vhd:4063:100  */
  assign n9133 = n9131 & n9132;
  /* TG68KdotC_Kernel.vhd:4063:83  */
  assign n9134 = n9129 | n9133;
  /* TG68KdotC_Kernel.vhd:4063:122  */
  assign n9135 = flags[2]; // extract
  /* TG68KdotC_Kernel.vhd:4063:114  */
  assign n9136 = n9134 | n9135;
  /* TG68KdotC_Kernel.vhd:4063:25  */
  assign n9138 = n9042 == 4'b1111;
  assign n9139 = {n9138, n9125, n9108, n9097, n9086, n9083, n9079, n9076, n9072, n9069, n9065, n9062, n9058, n9053, n9046, n9044};
  /* TG68KdotC_Kernel.vhd:4047:17  */
  always @*
    case (n9139)
      16'b1000000000000000: n9142 = n9136;
      16'b0100000000000000: n9142 = n9123;
      16'b0010000000000000: n9142 = n9106;
      16'b0001000000000000: n9142 = n9095;
      16'b0000100000000000: n9142 = n9084;
      16'b0000010000000000: n9142 = n9081;
      16'b0000001000000000: n9142 = n9077;
      16'b0000000100000000: n9142 = n9074;
      16'b0000000010000000: n9142 = n9070;
      16'b0000000001000000: n9142 = n9067;
      16'b0000000000100000: n9142 = n9063;
      16'b0000000000010000: n9142 = n9060;
      16'b0000000000001000: n9142 = n9056;
      16'b0000000000000100: n9142 = n9051;
      16'b0000000000000010: n9142 = 1'b0;
      16'b0000000000000001: n9142 = 1'b1;
      default: n9142 = exe_condition;
    endcase
  /* TG68KdotC_Kernel.vhd:4075:54  */
  assign n9147 = exec[69]; // extract
  /* TG68KdotC_Kernel.vhd:4077:60  */
  assign n9148 = data_read[15:0]; // extract
  /* TG68KdotC_Kernel.vhd:4078:43  */
  assign n9149 = exec[69]; // extract
  /* TG68KdotC_Kernel.vhd:4078:68  */
  assign n9150 = set[69]; // extract
  /* TG68KdotC_Kernel.vhd:4078:62  */
  assign n9151 = n9149 | n9150;
  /* TG68KdotC_Kernel.vhd:4080:49  */
  assign n9154 = movem_regaddr == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4081:49  */
  assign n9157 = movem_regaddr == 4'b0001;
  /* TG68KdotC_Kernel.vhd:4082:49  */
  assign n9160 = movem_regaddr == 4'b0010;
  /* TG68KdotC_Kernel.vhd:4083:49  */
  assign n9163 = movem_regaddr == 4'b0011;
  /* TG68KdotC_Kernel.vhd:4084:49  */
  assign n9166 = movem_regaddr == 4'b0100;
  /* TG68KdotC_Kernel.vhd:4085:49  */
  assign n9169 = movem_regaddr == 4'b0101;
  /* TG68KdotC_Kernel.vhd:4086:49  */
  assign n9172 = movem_regaddr == 4'b0110;
  /* TG68KdotC_Kernel.vhd:4087:49  */
  assign n9175 = movem_regaddr == 4'b0111;
  /* TG68KdotC_Kernel.vhd:4088:49  */
  assign n9178 = movem_regaddr == 4'b1000;
  /* TG68KdotC_Kernel.vhd:4089:49  */
  assign n9181 = movem_regaddr == 4'b1001;
  /* TG68KdotC_Kernel.vhd:4090:49  */
  assign n9184 = movem_regaddr == 4'b1010;
  /* TG68KdotC_Kernel.vhd:4091:49  */
  assign n9187 = movem_regaddr == 4'b1011;
  /* TG68KdotC_Kernel.vhd:4092:49  */
  assign n9190 = movem_regaddr == 4'b1100;
  /* TG68KdotC_Kernel.vhd:4093:49  */
  assign n9193 = movem_regaddr == 4'b1101;
  /* TG68KdotC_Kernel.vhd:4094:49  */
  assign n9196 = movem_regaddr == 4'b1110;
  /* TG68KdotC_Kernel.vhd:4095:49  */
  assign n9199 = movem_regaddr == 4'b1111;
  assign n9200 = {n9199, n9196, n9193, n9190, n9187, n9184, n9181, n9178, n9175, n9172, n9169, n9166, n9163, n9160, n9157, n9154};
  assign n9201 = sndopc[0]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9202 = n9201;
      16'b0100000000000000: n9202 = n9201;
      16'b0010000000000000: n9202 = n9201;
      16'b0001000000000000: n9202 = n9201;
      16'b0000100000000000: n9202 = n9201;
      16'b0000010000000000: n9202 = n9201;
      16'b0000001000000000: n9202 = n9201;
      16'b0000000100000000: n9202 = n9201;
      16'b0000000010000000: n9202 = n9201;
      16'b0000000001000000: n9202 = n9201;
      16'b0000000000100000: n9202 = n9201;
      16'b0000000000010000: n9202 = n9201;
      16'b0000000000001000: n9202 = n9201;
      16'b0000000000000100: n9202 = n9201;
      16'b0000000000000010: n9202 = n9201;
      16'b0000000000000001: n9202 = 1'b0;
      default: n9202 = n9201;
    endcase
  assign n9203 = sndopc[1]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9204 = n9203;
      16'b0100000000000000: n9204 = n9203;
      16'b0010000000000000: n9204 = n9203;
      16'b0001000000000000: n9204 = n9203;
      16'b0000100000000000: n9204 = n9203;
      16'b0000010000000000: n9204 = n9203;
      16'b0000001000000000: n9204 = n9203;
      16'b0000000100000000: n9204 = n9203;
      16'b0000000010000000: n9204 = n9203;
      16'b0000000001000000: n9204 = n9203;
      16'b0000000000100000: n9204 = n9203;
      16'b0000000000010000: n9204 = n9203;
      16'b0000000000001000: n9204 = n9203;
      16'b0000000000000100: n9204 = n9203;
      16'b0000000000000010: n9204 = 1'b0;
      16'b0000000000000001: n9204 = n9203;
      default: n9204 = n9203;
    endcase
  assign n9205 = sndopc[2]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9206 = n9205;
      16'b0100000000000000: n9206 = n9205;
      16'b0010000000000000: n9206 = n9205;
      16'b0001000000000000: n9206 = n9205;
      16'b0000100000000000: n9206 = n9205;
      16'b0000010000000000: n9206 = n9205;
      16'b0000001000000000: n9206 = n9205;
      16'b0000000100000000: n9206 = n9205;
      16'b0000000010000000: n9206 = n9205;
      16'b0000000001000000: n9206 = n9205;
      16'b0000000000100000: n9206 = n9205;
      16'b0000000000010000: n9206 = n9205;
      16'b0000000000001000: n9206 = n9205;
      16'b0000000000000100: n9206 = 1'b0;
      16'b0000000000000010: n9206 = n9205;
      16'b0000000000000001: n9206 = n9205;
      default: n9206 = n9205;
    endcase
  assign n9207 = sndopc[3]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9208 = n9207;
      16'b0100000000000000: n9208 = n9207;
      16'b0010000000000000: n9208 = n9207;
      16'b0001000000000000: n9208 = n9207;
      16'b0000100000000000: n9208 = n9207;
      16'b0000010000000000: n9208 = n9207;
      16'b0000001000000000: n9208 = n9207;
      16'b0000000100000000: n9208 = n9207;
      16'b0000000010000000: n9208 = n9207;
      16'b0000000001000000: n9208 = n9207;
      16'b0000000000100000: n9208 = n9207;
      16'b0000000000010000: n9208 = n9207;
      16'b0000000000001000: n9208 = 1'b0;
      16'b0000000000000100: n9208 = n9207;
      16'b0000000000000010: n9208 = n9207;
      16'b0000000000000001: n9208 = n9207;
      default: n9208 = n9207;
    endcase
  assign n9209 = sndopc[4]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9210 = n9209;
      16'b0100000000000000: n9210 = n9209;
      16'b0010000000000000: n9210 = n9209;
      16'b0001000000000000: n9210 = n9209;
      16'b0000100000000000: n9210 = n9209;
      16'b0000010000000000: n9210 = n9209;
      16'b0000001000000000: n9210 = n9209;
      16'b0000000100000000: n9210 = n9209;
      16'b0000000010000000: n9210 = n9209;
      16'b0000000001000000: n9210 = n9209;
      16'b0000000000100000: n9210 = n9209;
      16'b0000000000010000: n9210 = 1'b0;
      16'b0000000000001000: n9210 = n9209;
      16'b0000000000000100: n9210 = n9209;
      16'b0000000000000010: n9210 = n9209;
      16'b0000000000000001: n9210 = n9209;
      default: n9210 = n9209;
    endcase
  assign n9211 = sndopc[5]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9212 = n9211;
      16'b0100000000000000: n9212 = n9211;
      16'b0010000000000000: n9212 = n9211;
      16'b0001000000000000: n9212 = n9211;
      16'b0000100000000000: n9212 = n9211;
      16'b0000010000000000: n9212 = n9211;
      16'b0000001000000000: n9212 = n9211;
      16'b0000000100000000: n9212 = n9211;
      16'b0000000010000000: n9212 = n9211;
      16'b0000000001000000: n9212 = n9211;
      16'b0000000000100000: n9212 = 1'b0;
      16'b0000000000010000: n9212 = n9211;
      16'b0000000000001000: n9212 = n9211;
      16'b0000000000000100: n9212 = n9211;
      16'b0000000000000010: n9212 = n9211;
      16'b0000000000000001: n9212 = n9211;
      default: n9212 = n9211;
    endcase
  assign n9213 = sndopc[6]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9214 = n9213;
      16'b0100000000000000: n9214 = n9213;
      16'b0010000000000000: n9214 = n9213;
      16'b0001000000000000: n9214 = n9213;
      16'b0000100000000000: n9214 = n9213;
      16'b0000010000000000: n9214 = n9213;
      16'b0000001000000000: n9214 = n9213;
      16'b0000000100000000: n9214 = n9213;
      16'b0000000010000000: n9214 = n9213;
      16'b0000000001000000: n9214 = 1'b0;
      16'b0000000000100000: n9214 = n9213;
      16'b0000000000010000: n9214 = n9213;
      16'b0000000000001000: n9214 = n9213;
      16'b0000000000000100: n9214 = n9213;
      16'b0000000000000010: n9214 = n9213;
      16'b0000000000000001: n9214 = n9213;
      default: n9214 = n9213;
    endcase
  assign n9215 = sndopc[7]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9216 = n9215;
      16'b0100000000000000: n9216 = n9215;
      16'b0010000000000000: n9216 = n9215;
      16'b0001000000000000: n9216 = n9215;
      16'b0000100000000000: n9216 = n9215;
      16'b0000010000000000: n9216 = n9215;
      16'b0000001000000000: n9216 = n9215;
      16'b0000000100000000: n9216 = n9215;
      16'b0000000010000000: n9216 = 1'b0;
      16'b0000000001000000: n9216 = n9215;
      16'b0000000000100000: n9216 = n9215;
      16'b0000000000010000: n9216 = n9215;
      16'b0000000000001000: n9216 = n9215;
      16'b0000000000000100: n9216 = n9215;
      16'b0000000000000010: n9216 = n9215;
      16'b0000000000000001: n9216 = n9215;
      default: n9216 = n9215;
    endcase
  assign n9217 = sndopc[8]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9218 = n9217;
      16'b0100000000000000: n9218 = n9217;
      16'b0010000000000000: n9218 = n9217;
      16'b0001000000000000: n9218 = n9217;
      16'b0000100000000000: n9218 = n9217;
      16'b0000010000000000: n9218 = n9217;
      16'b0000001000000000: n9218 = n9217;
      16'b0000000100000000: n9218 = 1'b0;
      16'b0000000010000000: n9218 = n9217;
      16'b0000000001000000: n9218 = n9217;
      16'b0000000000100000: n9218 = n9217;
      16'b0000000000010000: n9218 = n9217;
      16'b0000000000001000: n9218 = n9217;
      16'b0000000000000100: n9218 = n9217;
      16'b0000000000000010: n9218 = n9217;
      16'b0000000000000001: n9218 = n9217;
      default: n9218 = n9217;
    endcase
  assign n9219 = sndopc[9]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9220 = n9219;
      16'b0100000000000000: n9220 = n9219;
      16'b0010000000000000: n9220 = n9219;
      16'b0001000000000000: n9220 = n9219;
      16'b0000100000000000: n9220 = n9219;
      16'b0000010000000000: n9220 = n9219;
      16'b0000001000000000: n9220 = 1'b0;
      16'b0000000100000000: n9220 = n9219;
      16'b0000000010000000: n9220 = n9219;
      16'b0000000001000000: n9220 = n9219;
      16'b0000000000100000: n9220 = n9219;
      16'b0000000000010000: n9220 = n9219;
      16'b0000000000001000: n9220 = n9219;
      16'b0000000000000100: n9220 = n9219;
      16'b0000000000000010: n9220 = n9219;
      16'b0000000000000001: n9220 = n9219;
      default: n9220 = n9219;
    endcase
  assign n9221 = sndopc[10]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9222 = n9221;
      16'b0100000000000000: n9222 = n9221;
      16'b0010000000000000: n9222 = n9221;
      16'b0001000000000000: n9222 = n9221;
      16'b0000100000000000: n9222 = n9221;
      16'b0000010000000000: n9222 = 1'b0;
      16'b0000001000000000: n9222 = n9221;
      16'b0000000100000000: n9222 = n9221;
      16'b0000000010000000: n9222 = n9221;
      16'b0000000001000000: n9222 = n9221;
      16'b0000000000100000: n9222 = n9221;
      16'b0000000000010000: n9222 = n9221;
      16'b0000000000001000: n9222 = n9221;
      16'b0000000000000100: n9222 = n9221;
      16'b0000000000000010: n9222 = n9221;
      16'b0000000000000001: n9222 = n9221;
      default: n9222 = n9221;
    endcase
  assign n9223 = sndopc[11]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9224 = n9223;
      16'b0100000000000000: n9224 = n9223;
      16'b0010000000000000: n9224 = n9223;
      16'b0001000000000000: n9224 = n9223;
      16'b0000100000000000: n9224 = 1'b0;
      16'b0000010000000000: n9224 = n9223;
      16'b0000001000000000: n9224 = n9223;
      16'b0000000100000000: n9224 = n9223;
      16'b0000000010000000: n9224 = n9223;
      16'b0000000001000000: n9224 = n9223;
      16'b0000000000100000: n9224 = n9223;
      16'b0000000000010000: n9224 = n9223;
      16'b0000000000001000: n9224 = n9223;
      16'b0000000000000100: n9224 = n9223;
      16'b0000000000000010: n9224 = n9223;
      16'b0000000000000001: n9224 = n9223;
      default: n9224 = n9223;
    endcase
  assign n9225 = sndopc[12]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9226 = n9225;
      16'b0100000000000000: n9226 = n9225;
      16'b0010000000000000: n9226 = n9225;
      16'b0001000000000000: n9226 = 1'b0;
      16'b0000100000000000: n9226 = n9225;
      16'b0000010000000000: n9226 = n9225;
      16'b0000001000000000: n9226 = n9225;
      16'b0000000100000000: n9226 = n9225;
      16'b0000000010000000: n9226 = n9225;
      16'b0000000001000000: n9226 = n9225;
      16'b0000000000100000: n9226 = n9225;
      16'b0000000000010000: n9226 = n9225;
      16'b0000000000001000: n9226 = n9225;
      16'b0000000000000100: n9226 = n9225;
      16'b0000000000000010: n9226 = n9225;
      16'b0000000000000001: n9226 = n9225;
      default: n9226 = n9225;
    endcase
  assign n9227 = sndopc[13]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9228 = n9227;
      16'b0100000000000000: n9228 = n9227;
      16'b0010000000000000: n9228 = 1'b0;
      16'b0001000000000000: n9228 = n9227;
      16'b0000100000000000: n9228 = n9227;
      16'b0000010000000000: n9228 = n9227;
      16'b0000001000000000: n9228 = n9227;
      16'b0000000100000000: n9228 = n9227;
      16'b0000000010000000: n9228 = n9227;
      16'b0000000001000000: n9228 = n9227;
      16'b0000000000100000: n9228 = n9227;
      16'b0000000000010000: n9228 = n9227;
      16'b0000000000001000: n9228 = n9227;
      16'b0000000000000100: n9228 = n9227;
      16'b0000000000000010: n9228 = n9227;
      16'b0000000000000001: n9228 = n9227;
      default: n9228 = n9227;
    endcase
  assign n9229 = sndopc[14]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9230 = n9229;
      16'b0100000000000000: n9230 = 1'b0;
      16'b0010000000000000: n9230 = n9229;
      16'b0001000000000000: n9230 = n9229;
      16'b0000100000000000: n9230 = n9229;
      16'b0000010000000000: n9230 = n9229;
      16'b0000001000000000: n9230 = n9229;
      16'b0000000100000000: n9230 = n9229;
      16'b0000000010000000: n9230 = n9229;
      16'b0000000001000000: n9230 = n9229;
      16'b0000000000100000: n9230 = n9229;
      16'b0000000000010000: n9230 = n9229;
      16'b0000000000001000: n9230 = n9229;
      16'b0000000000000100: n9230 = n9229;
      16'b0000000000000010: n9230 = n9229;
      16'b0000000000000001: n9230 = n9229;
      default: n9230 = n9229;
    endcase
  assign n9231 = sndopc[15]; // extract
  /* TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9200)
      16'b1000000000000000: n9232 = 1'b0;
      16'b0100000000000000: n9232 = n9231;
      16'b0010000000000000: n9232 = n9231;
      16'b0001000000000000: n9232 = n9231;
      16'b0000100000000000: n9232 = n9231;
      16'b0000010000000000: n9232 = n9231;
      16'b0000001000000000: n9232 = n9231;
      16'b0000000100000000: n9232 = n9231;
      16'b0000000010000000: n9232 = n9231;
      16'b0000000001000000: n9232 = n9231;
      16'b0000000000100000: n9232 = n9231;
      16'b0000000000010000: n9232 = n9231;
      16'b0000000000001000: n9232 = n9231;
      16'b0000000000000100: n9232 = n9231;
      16'b0000000000000010: n9232 = n9231;
      16'b0000000000000001: n9232 = n9231;
      default: n9232 = n9231;
    endcase
  assign n9233 = {n9232, n9230, n9228, n9226, n9224, n9222, n9220, n9218, n9216, n9214, n9212, n9210, n9208, n9206, n9204, n9202};
  /* TG68KdotC_Kernel.vhd:4078:33  */
  assign n9234 = n9151 ? n9233 : sndopc;
  /* TG68KdotC_Kernel.vhd:4076:33  */
  assign n9235 = decodeopc ? n9148 : n9234;
  /* TG68KdotC_Kernel.vhd:4107:26  */
  assign n9243 = sndopc[3:0]; // extract
  /* TG68KdotC_Kernel.vhd:4107:38  */
  assign n9245 = n9243 == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4108:34  */
  assign n9246 = sndopc[7:4]; // extract
  /* TG68KdotC_Kernel.vhd:4108:46  */
  assign n9248 = n9246 == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4110:42  */
  assign n9250 = sndopc[11:8]; // extract
  /* TG68KdotC_Kernel.vhd:4110:55  */
  assign n9252 = n9250 == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4111:50  */
  assign n9253 = sndopc[15:12]; // extract
  /* TG68KdotC_Kernel.vhd:4111:64  */
  assign n9255 = n9253 == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4111:41  */
  assign n9258 = n9255 ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:4115:60  */
  assign n9260 = sndopc[15:12]; // extract
  /* TG68KdotC_Kernel.vhd:4117:60  */
  assign n9261 = sndopc[11:8]; // extract
  /* TG68KdotC_Kernel.vhd:4110:33  */
  assign n9263 = n9252 ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:4110:33  */
  assign n9264 = n9252 ? n9260 : n9261;
  /* TG68KdotC_Kernel.vhd:4110:33  */
  assign n9266 = n9252 ? n9258 : 1'b1;
  /* TG68KdotC_Kernel.vhd:4120:52  */
  assign n9267 = sndopc[7:4]; // extract
  assign n9269 = {1'b1, n9263};
  assign n9270 = n9269[0]; // extract
  /* TG68KdotC_Kernel.vhd:4108:25  */
  assign n9271 = n9248 ? n9270 : 1'b1;
  assign n9272 = n9269[1]; // extract
  /* TG68KdotC_Kernel.vhd:4108:25  */
  assign n9274 = n9248 ? n9272 : 1'b0;
  /* TG68KdotC_Kernel.vhd:4108:25  */
  assign n9275 = n9248 ? n9264 : n9267;
  /* TG68KdotC_Kernel.vhd:4108:25  */
  assign n9277 = n9248 ? n9266 : 1'b1;
  /* TG68KdotC_Kernel.vhd:4124:44  */
  assign n9278 = sndopc[3:0]; // extract
  assign n9279 = {n9274, n9271};
  /* TG68KdotC_Kernel.vhd:4107:17  */
  assign n9281 = n9245 ? n9279 : 2'b00;
  /* TG68KdotC_Kernel.vhd:4107:17  */
  assign n9284 = n9245 ? n9275 : n9278;
  /* TG68KdotC_Kernel.vhd:4107:17  */
  assign n9286 = n9245 ? n9277 : 1'b1;
  /* TG68KdotC_Kernel.vhd:4126:29  */
  assign n9288 = movem_mux[1:0]; // extract
  /* TG68KdotC_Kernel.vhd:4126:41  */
  assign n9290 = n9288 == 2'b00;
  /* TG68KdotC_Kernel.vhd:4128:37  */
  assign n9292 = movem_mux[2]; // extract
  /* TG68KdotC_Kernel.vhd:4128:40  */
  assign n9293 = ~n9292;
  assign n9295 = n9282[0]; // extract
  /* TG68KdotC_Kernel.vhd:4128:25  */
  assign n9296 = n9293 ? 1'b1 : n9295;
  /* TG68KdotC_Kernel.vhd:4132:37  */
  assign n9297 = movem_mux[0]; // extract
  /* TG68KdotC_Kernel.vhd:4132:40  */
  assign n9298 = ~n9297;
  assign n9300 = n9282[0]; // extract
  /* TG68KdotC_Kernel.vhd:4132:25  */
  assign n9301 = n9298 ? 1'b1 : n9300;
  assign n9302 = {1'b1, n9296};
  assign n9303 = n9302[0]; // extract
  /* TG68KdotC_Kernel.vhd:4126:17  */
  assign n9304 = n9290 ? n9303 : n9301;
  assign n9305 = n9302[1]; // extract
  assign n9306 = n9282[1]; // extract
  /* TG68KdotC_Kernel.vhd:4126:17  */
  assign n9307 = n9290 ? n9305 : n9306;
  /* TG68KdotC_Kernel.vhd:464:17  */
  always @(posedge clk)
    n9310 <= n106;
  /* TG68KdotC_Kernel.vhd:458:17  */
  assign n9311 = clkena_in ? n87 : syncreset;
  /* TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n83)
    if (n83)
      n9312 <= 4'b0000;
    else
      n9312 <= n9311;
  /* TG68KdotC_Kernel.vhd:458:17  */
  assign n9313 = clkena_in ? n89 : reset;
  /* TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n83)
    if (n83)
      n9314 <= 1'b1;
    else
      n9314 <= n9313;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9315 <= n1423;
  /* TG68KdotC_Kernel.vhd:941:17  */
  assign n9316 = n983 ? addr : tmp_tg68_pc;
  /* TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9317 <= n9316;
  /* TG68KdotC_Kernel.vhd:941:17  */
  assign n9318 = n984 ? addr : memaddr;
  /* TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9319 <= n9318;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9320 <= n1425;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9321 <= n1426;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9322 <= n1428;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9323 <= n1430;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9324 <= n1431;
  /* TG68KdotC_Kernel.vhd:4073:17  */
  assign n9325 = clkena_lw ? n9235 : sndopc;
  /* TG68KdotC_Kernel.vhd:4073:17  */
  always @(posedge clk)
    n9326 <= n9325;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9327 <= n1432;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9328 <= n1433;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9329 <= n1435;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9331 = clkena_lw ? rf_source_addr : rf_source_addrd;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9332 <= n9331;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9333 = {n309, n304, n306};
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9336 = clkena_lw ? rf_dest_addr : rdindex_a;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9337 <= n9336;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9338 = clkena_lw ? rf_source_addr : rdindex_b;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9339 <= n9338;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9340 = clkena_lw ? n268 : wr_areg;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9341 <= n9340;
  /* TG68KdotC_Kernel.vhd:941:17  */
  assign n9342 = clkena_in ? n970 : memaddr_delta_rega;
  /* TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9343 <= n9342;
  /* TG68KdotC_Kernel.vhd:941:17  */
  assign n9344 = clkena_in ? n972 : memaddr_delta_regb;
  /* TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9345 <= n9344;
  /* TG68KdotC_Kernel.vhd:941:17  */
  assign n9346 = clkena_in ? n975 : use_base;
  /* TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9347 <= n9346;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9348 <= n711;
  /* TG68KdotC_Kernel.vhd:743:9  */
  assign n9349 = {n566, n567};
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9351 <= n712;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9352 <= n1436;
  assign n9354 = {n908, n905};
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9355 <= n1438;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9356 <= n1439;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9357 <= n714;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9358 <= n1441;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9359 <= n1443;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9360 <= n716;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9361 <= n1445;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9362 <= n1447;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9363 <= n1449;
  /* TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9364 <= n1763;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9365 <= n717;
  /* TG68KdotC_Kernel.vhd:1254:17  */
  assign n9366 = clkena_lw ? n1558 : exec_tas;
  /* TG68KdotC_Kernel.vhd:1254:17  */
  always @(posedge clk)
    n9367 <= n9366;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9368 <= n1450;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9369 <= n1452;
  /* TG68KdotC_Kernel.vhd:4073:17  */
  assign n9370 = clkena_lw ? n9147 : movem_actiond;
  /* TG68KdotC_Kernel.vhd:4073:17  */
  always @(posedge clk)
    n9371 <= n9370;
  /* TG68KdotC_Kernel.vhd:4073:17  */
  assign n9372 = {n9281, n9307, n9304};
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9374 <= n719;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9375 <= n721;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9376 <= n1454;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9377 <= n1456;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9378 <= n1458;
  /* TG68KdotC_Kernel.vhd:3239:17  */
  always @(posedge clk)
    n9379 <= n7844;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9380 <= n1459;
  /* TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9381 <= n1765;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9382 <= n1461;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9383 <= n722;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9384 <= n1463;
  /* TG68KdotC_Kernel.vhd:870:17  */
  assign n9385 = clkena_lw ? n834 : trap_vector;
  /* TG68KdotC_Kernel.vhd:870:17  */
  always @(posedge clk)
    n9386 <= n9385;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9387 = n283 ? reg_qa : usp;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9388 <= n9387;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9389 <= n1464;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9390 <= n1465;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9391 <= n1467;
  /* TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9392 <= n1767;
  /* TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9393 <= n1769;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9394 <= n1469;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9395 <= n724;
  /* TG68KdotC_Kernel.vhd:743:9  */
  assign n9396 = {n148, n149};
  /* TG68KdotC_Kernel.vhd:484:17  */
  assign n9397 = n153 ? n158 : bf_ext_in;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9398 <= n9397;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9399 <= n1471;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9400 <= n1472;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9401 <= n1473;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9402 <= n1474;
  /* TG68KdotC_Kernel.vhd:1254:17  */
  always @(posedge clk)
    n9403 <= n1528;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9404 <= n205;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9405 <= n206;
  /* TG68KdotC_Kernel.vhd:484:17  */
  assign n9406 = {n1643, n1642, n1644};
  assign n9407 = {1'b0, n1598};
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9408 <= n1475;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9409 <= n1476;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  assign n9410 = {1'b0, n1609};
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9411 <= n1477;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9412 <= n1478;
  /* TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9413 <= n9009;
  /* TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9414 <= n9011;
  /* TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9415 <= n9012;
  /* TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9416 <= n9013;
  /* TG68KdotC_Kernel.vhd:4008:9  */
  assign n9417 = {n8918, n8916, n8914, n8913, n8912, n8911, n8910, n7647, n7606, n8909, n8925, n7604, n8907, n8906, n7599, n8905, n8904, n8903, n8902, n8924, n8900, n8923, n8898, n7592, n8921, n8897, n8895, n8893, n8892, n7581, n7578, n7575, n8891, n8890, n7567, n8889, n8888, n8887, n7556, n7554, n7551, n1879, n8886, n8885, n8884, n8883, n7541, n8882, n8881, n7624, n7537, n8919, n8880, n8878, n8877, n8876, n7619, n8875, n8874, n8873, n7529, n7617, n8872};
  assign n9418 = {n7720, n7757, n7718, n7756, n7716, n7714, n7753, n7712, n7751, n7833, n7708, n7706, n7704, n7746, n7832, n7744, n7831, n8929, n8928, n8930, n7698, n7740, n7696, n7694, n7692, n7690, n7688, n7686, n7684, n7682, n7680, n7677, n7673, n7669, n7666, n7663, n7659, n7656, n7653};
  /* TG68KdotC_Kernel.vhd:1254:17  */
  assign n9419 = clkena_lw ? n1568 : exec;
  /* TG68KdotC_Kernel.vhd:1254:17  */
  always @(posedge clk)
    n9420 <= n9419;
  /* TG68KdotC_Kernel.vhd:3239:17  */
  always @(posedge clk)
    n9421 <= n7846;
  /* TG68KdotC_Kernel.vhd:3239:17  */
  assign n9422 = {n255, n254};
  /* TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9423 <= n1761;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9424 <= n1421;
  /* TG68KdotC_Kernel.vhd:1053:17  */
  assign n9425 = {n9423, n9424};
  /* TG68KdotC_Kernel.vhd:559:35  */
  reg [31:0] regfile[15:0] ; // memory
  initial begin
    regfile[15] = 32'b00000000000000000000000000000000;
    regfile[14] = 32'b00000000000000000000000000000000;
    regfile[13] = 32'b00000000000000000000000000000000;
    regfile[12] = 32'b00000000000000000000000000000000;
    regfile[11] = 32'b00000000000000000000000000000000;
    regfile[10] = 32'b00000000000000000000000000000000;
    regfile[9] = 32'b00000000000000000000000000000000;
    regfile[8] = 32'b00000000000000000000000000000000;
    regfile[7] = 32'b00000000000000000000000000000000;
    regfile[6] = 32'b00000000000000000000000000000000;
    regfile[5] = 32'b00000000000000000000000000000000;
    regfile[4] = 32'b00000000000000000000000000000000;
    regfile[3] = 32'b00000000000000000000000000000000;
    regfile[2] = 32'b00000000000000000000000000000000;
    regfile[1] = 32'b00000000000000000000000000000000;
    regfile[0] = 32'b00000000000000000000000000000000;
    end
  assign n9428 = regfile[rdindex_b];
  assign n9429 = regfile[rdindex_a];
  always @(posedge clk)
    if (n279)
      regfile[rdindex_a] <= regin;
  /* TG68KdotC_Kernel.vhd:559:35  */
  /* TG68KdotC_Kernel.vhd:558:35  */
  /* TG68KdotC_Kernel.vhd:567:49  */
endmodule

