module tg68k_fpu_packeddecimal
  (input  clk,
   input  nreset,
   input  clkena,
   input  start_conversion,
   input  packed_to_extended,
   input  [6:0] k_factor,
   input  [79:0] extended_in,
   input  [95:0] packed_in,
   output conversion_done,
   output conversion_valid,
   output [79:0] extended_out,
   output [95:0] packed_out,
   output overflow,
   output inexact,
   output invalid);
  reg [2:0] packed_state;
  wire [67:0] bcd_digits;
  wire [11:0] bcd_exponent;
  wire [63:0] binary_mantissa;
  wire [10:0] decimal_exponent;
  wire [127:0] work_mantissa;
  wire [31:0] work_exponent;
  wire result_sign;
  wire exp_sign;
  wire [5:0] cycle_count;
  reg [127:0] packed_conversion_temp_mantissa;
  wire n15692;
  wire [2:0] n15695;
  wire n15697;
  wire n15698;
  wire n15699;
  wire [11:0] n15700;
  wire [67:0] n15701;
  wire [3:0] n15702;
  wire n15704;
  wire n15707;
  wire [3:0] n15709;
  wire n15711;
  wire n15713;
  wire [3:0] n15714;
  wire n15716;
  wire n15718;
  wire [3:0] n15719;
  wire n15721;
  wire n15723;
  wire [3:0] n15724;
  wire n15726;
  wire n15728;
  wire [3:0] n15729;
  wire n15731;
  wire n15733;
  wire [3:0] n15734;
  wire n15736;
  wire n15738;
  wire [3:0] n15739;
  wire n15741;
  wire n15743;
  wire [3:0] n15744;
  wire n15746;
  wire n15748;
  wire [3:0] n15749;
  wire n15751;
  wire n15753;
  wire [3:0] n15754;
  wire n15756;
  wire n15758;
  wire [3:0] n15759;
  wire n15761;
  wire n15763;
  wire [3:0] n15764;
  wire n15766;
  wire n15768;
  wire [3:0] n15769;
  wire n15771;
  wire n15773;
  wire [3:0] n15774;
  wire n15776;
  wire n15778;
  wire [3:0] n15779;
  wire n15781;
  wire n15783;
  wire [3:0] n15784;
  wire n15786;
  wire n15788;
  wire [3:0] n15789;
  wire n15791;
  wire n15793;
  wire [3:0] n15794;
  wire n15796;
  wire n15798;
  wire [3:0] n15799;
  wire n15801;
  wire n15803;
  wire n15804;
  wire [14:0] n15805;
  wire [30:0] n15806;
  wire [31:0] n15807;
  wire [31:0] n15809;
  wire [63:0] n15810;
  wire [14:0] n15812;
  wire n15814;
  wire n15815;
  wire [62:0] n15816;
  wire n15818;
  wire n15819;
  wire [95:0] n15838;
  wire n15840;
  wire n15842;
  wire [2:0] n15844;
  wire [67:0] n15845;
  wire [67:0] n15846;
  wire [11:0] n15848;
  wire [78:0] n15849;
  wire n15851;
  wire [95:0] n15853;
  wire [2:0] n15856;
  wire [95:0] n15857;
  wire n15858;
  wire n15859;
  wire [2:0] n15860;
  wire n15861;
  wire n15862;
  wire [95:0] n15863;
  wire n15864;
  wire n15865;
  wire [2:0] n15867;
  wire [67:0] n15868;
  wire [11:0] n15869;
  wire [127:0] n15870;
  wire [127:0] n15871;
  wire [31:0] n15872;
  wire n15873;
  wire n15874;
  wire n15876;
  wire [31:0] n15877;
  wire n15879;
  wire [63:0] n15881;
  wire [127:0] n15883;
  wire [31:0] n15884;
  wire n15886;
  wire [3:0] n15887;
  wire [30:0] n15888;
  wire [31:0] n15889;
  wire n15891;
  wire [3:0] n15892;
  wire [30:0] n15893;
  wire [31:0] n15894;
  wire n15896;
  wire [3:0] n15897;
  wire [30:0] n15898;
  wire [31:0] n15899;
  wire n15901;
  wire [3:0] n15902;
  wire [30:0] n15903;
  wire [31:0] n15904;
  wire n15906;
  wire [3:0] n15907;
  wire [30:0] n15908;
  wire [31:0] n15909;
  wire n15911;
  wire [3:0] n15912;
  wire [30:0] n15913;
  wire [31:0] n15914;
  wire n15916;
  wire [3:0] n15917;
  wire [30:0] n15918;
  wire [31:0] n15919;
  wire n15921;
  wire [3:0] n15922;
  wire [30:0] n15923;
  wire [31:0] n15924;
  wire n15926;
  wire [3:0] n15927;
  wire [30:0] n15928;
  wire [31:0] n15929;
  wire n15931;
  wire [3:0] n15932;
  wire [30:0] n15933;
  wire [31:0] n15934;
  wire n15936;
  wire [3:0] n15937;
  wire [30:0] n15938;
  wire [31:0] n15939;
  wire n15941;
  wire [3:0] n15942;
  wire [30:0] n15943;
  wire [31:0] n15944;
  wire n15946;
  wire [3:0] n15947;
  wire [30:0] n15948;
  wire [31:0] n15949;
  wire n15951;
  wire [3:0] n15952;
  wire [30:0] n15953;
  wire [31:0] n15954;
  wire n15956;
  wire [3:0] n15957;
  wire [30:0] n15958;
  wire [31:0] n15959;
  wire n15961;
  wire [3:0] n15962;
  wire [30:0] n15963;
  wire [31:0] n15964;
  wire n15966;
  wire [3:0] n15967;
  wire [30:0] n15968;
  wire [31:0] n15969;
  wire n15971;
  wire [16:0] n15972;
  reg [31:0] n15974;
  wire [255:0] n15975;
  wire [255:0] n15977;
  wire [127:0] n15978;
  wire [30:0] n15979;
  wire [127:0] n15980;
  wire [127:0] n15981;
  wire [31:0] n15982;
  wire [31:0] n15984;
  wire [5:0] n15985;
  wire [3:0] n15994;
  wire [30:0] n15995;
  wire [31:0] n15996;
  wire [3:0] n15998;
  wire [30:0] n15999;
  wire [31:0] n16000;
  wire [3:0] n16002;
  wire [30:0] n16003;
  wire [31:0] n16004;
  wire n16007;
  wire n16009;
  wire n16010;
  wire n16012;
  wire n16013;
  wire n16017;
  wire [31:0] n16023;
  wire [31:0] n16025;
  wire [31:0] n16027;
  wire [31:0] n16028;
  wire [31:0] n16029;
  wire [31:0] n16034;
  wire [31:0] n16035;
  wire [31:0] n16036;
  wire [31:0] n16037;
  wire [10:0] n16038;
  wire [3:0] n16047;
  wire [30:0] n16048;
  wire [31:0] n16049;
  wire [3:0] n16051;
  wire [30:0] n16052;
  wire [31:0] n16053;
  wire [3:0] n16055;
  wire [30:0] n16056;
  wire [31:0] n16057;
  wire n16060;
  wire n16062;
  wire n16063;
  wire n16065;
  wire n16066;
  wire n16070;
  wire [31:0] n16076;
  wire [31:0] n16078;
  wire [31:0] n16080;
  wire [31:0] n16081;
  wire [31:0] n16082;
  wire [31:0] n16087;
  wire [31:0] n16088;
  wire [31:0] n16089;
  wire [10:0] n16090;
  wire [10:0] n16091;
  wire [63:0] n16092;
  wire [2:0] n16094;
  wire [63:0] n16095;
  wire [10:0] n16096;
  wire [5:0] n16098;
  wire [127:0] n16099;
  wire n16102;
  wire [31:0] n16103;
  wire n16105;
  wire n16107;
  wire [31:0] n16109;
  wire [31:0] n16111;
  wire [10:0] n16112;
  wire [31:0] n16114;
  wire [31:0] n16116;
  wire [31:0] n16117;
  wire [10:0] n16118;
  wire [10:0] n16119;
  wire n16122;
  wire [67:0] n16124;
  wire [10:0] n16125;
  wire n16126;
  wire [127:0] n16127;
  wire [31:0] n16128;
  wire n16130;
  wire [3:0] n16131;
  wire [3:0] n16133;
  wire n16135;
  wire [3:0] n16136;
  wire [3:0] n16138;
  wire n16140;
  wire [3:0] n16141;
  wire [3:0] n16143;
  wire n16145;
  wire [3:0] n16146;
  wire [3:0] n16148;
  wire n16150;
  wire [3:0] n16151;
  wire [3:0] n16153;
  wire n16155;
  wire [3:0] n16156;
  wire [3:0] n16158;
  wire n16160;
  wire [3:0] n16161;
  wire [3:0] n16163;
  wire n16165;
  wire [3:0] n16166;
  wire [3:0] n16168;
  wire n16170;
  wire [3:0] n16171;
  wire [3:0] n16173;
  wire n16175;
  wire [3:0] n16176;
  wire [3:0] n16178;
  wire n16180;
  wire [3:0] n16181;
  wire [3:0] n16183;
  wire n16185;
  wire [3:0] n16186;
  wire [3:0] n16188;
  wire n16190;
  wire [3:0] n16191;
  wire [3:0] n16193;
  wire n16195;
  wire [3:0] n16196;
  wire [3:0] n16198;
  wire n16200;
  wire [3:0] n16201;
  wire [3:0] n16203;
  wire n16205;
  wire [3:0] n16206;
  wire [3:0] n16208;
  wire n16210;
  wire [3:0] n16211;
  wire [3:0] n16213;
  wire n16215;
  wire [16:0] n16216;
  wire [3:0] n16217;
  reg [3:0] n16218;
  wire [3:0] n16219;
  reg [3:0] n16220;
  wire [3:0] n16221;
  reg [3:0] n16222;
  wire [3:0] n16223;
  reg [3:0] n16224;
  wire [3:0] n16225;
  reg [3:0] n16226;
  wire [3:0] n16227;
  reg [3:0] n16228;
  wire [3:0] n16229;
  reg [3:0] n16230;
  wire [3:0] n16231;
  reg [3:0] n16232;
  wire [3:0] n16233;
  reg [3:0] n16234;
  wire [3:0] n16235;
  reg [3:0] n16236;
  wire [3:0] n16237;
  reg [3:0] n16238;
  wire [3:0] n16239;
  reg [3:0] n16240;
  wire [3:0] n16241;
  reg [3:0] n16242;
  wire [3:0] n16243;
  reg [3:0] n16244;
  wire [3:0] n16245;
  reg [3:0] n16246;
  wire [3:0] n16247;
  reg [3:0] n16248;
  wire [3:0] n16249;
  reg [3:0] n16250;
  wire [31:0] n16251;
  wire [31:0] n16253;
  wire [5:0] n16254;
  wire [31:0] n16255;
  wire [31:0] n16256;
  wire [31:0] n16257;
  wire [10:0] n16258;
  wire [31:0] n16259;
  wire n16261;
  wire [31:0] n16263;
  wire [31:0] n16264;
  wire [31:0] n16271;
  wire [30:0] n16272;
  wire [3:0] n16273;
  wire [31:0] n16277;
  wire [31:0] n16279;
  wire [30:0] n16280;
  wire [3:0] n16281;
  wire [31:0] n16284;
  wire [31:0] n16286;
  wire [30:0] n16287;
  wire [3:0] n16288;
  wire [11:0] n16289;
  wire [31:0] n16291;
  wire [31:0] n16298;
  wire [30:0] n16299;
  wire [3:0] n16300;
  wire [31:0] n16304;
  wire [31:0] n16306;
  wire [30:0] n16307;
  wire [3:0] n16308;
  wire [31:0] n16311;
  wire [31:0] n16313;
  wire [30:0] n16314;
  wire [3:0] n16315;
  wire [11:0] n16316;
  wire [11:0] n16317;
  wire n16320;
  wire n16322;
  wire [2:0] n16324;
  wire [67:0] n16325;
  wire [67:0] n16326;
  wire [11:0] n16327;
  wire [10:0] n16328;
  wire n16329;
  wire [5:0] n16330;
  wire n16332;
  wire n16334;
  wire [31:0] n16335;
  wire [31:0] n16337;
  wire [31:0] n16339;
  wire [31:0] n16341;
  wire n16343;
  wire [79:0] n16345;
  wire n16347;
  wire [15:0] n16349;
  wire [16:0] n16351;
  wire [79:0] n16353;
  wire [30:0] n16354;
  wire [14:0] n16355;
  wire [15:0] n16356;
  wire [79:0] n16357;
  wire [79:0] n16358;
  wire n16360;
  wire [79:0] n16361;
  wire n16362;
  wire [79:0] n16364;
  wire n16365;
  wire n16368;
  wire n16370;
  wire n16371;
  wire [1:0] n16372;
  wire [3:0] n16374;
  wire [15:0] n16375;
  wire [16:0] n16377;
  wire [27:0] n16379;
  wire [95:0] n16380;
  wire [95:0] n16381;
  wire n16383;
  wire [6:0] n16384;
  reg n16388;
  reg n16392;
  reg [79:0] n16394;
  reg [95:0] n16396;
  reg n16399;
  reg n16403;
  reg n16406;
  reg [2:0] n16411;
  reg [67:0] n16413;
  reg [11:0] n16415;
  reg [63:0] n16417;
  reg [10:0] n16419;
  reg [127:0] n16421;
  reg [31:0] n16423;
  reg n16425;
  reg n16427;
  reg [5:0] n16430;
  reg [127:0] n16432;
  wire n16507;
  wire n16508;
  wire [127:0] n16509;
  reg [127:0] n16510;
  wire [2:0] n16519;
  reg [2:0] n16520;
  wire n16521;
  wire n16522;
  wire [67:0] n16523;
  reg [67:0] n16524;
  wire n16525;
  wire n16526;
  wire [11:0] n16527;
  reg [11:0] n16528;
  wire n16529;
  wire n16530;
  wire [63:0] n16531;
  reg [63:0] n16532;
  wire n16534;
  wire n16535;
  wire [10:0] n16536;
  reg [10:0] n16537;
  wire n16538;
  wire n16539;
  wire [127:0] n16540;
  reg [127:0] n16541;
  wire n16542;
  wire n16543;
  wire [31:0] n16544;
  reg [31:0] n16545;
  wire n16546;
  wire n16547;
  wire n16548;
  reg n16549;
  wire n16550;
  wire n16551;
  wire n16552;
  reg n16553;
  wire [5:0] n16554;
  reg [5:0] n16555;
  wire n16556;
  reg n16557;
  wire n16558;
  reg n16559;
  wire [79:0] n16560;
  reg [79:0] n16561;
  wire [95:0] n16562;
  reg [95:0] n16563;
  wire n16564;
  reg n16565;
  wire n16566;
  reg n16567;
  wire n16568;
  reg n16569;
  assign conversion_done = n16557; //(module output)
  assign conversion_valid = n16559; //(module output)
  assign extended_out = n16561; //(module output)
  assign packed_out = n16563; //(module output)
  assign overflow = n16565; //(module output)
  assign inexact = n16567; //(module output)
  assign invalid = n16569; //(module output)
  /* TG68K_FPU_PackedDecimal.vhd:78:12  */
  always @*
    packed_state = n16520; // (isignal)
  initial
    packed_state = 3'b000;
  /* TG68K_FPU_PackedDecimal.vhd:85:12  */
  assign bcd_digits = n16524; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:86:12  */
  assign bcd_exponent = n16528; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:87:12  */
  assign binary_mantissa = n16532; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:89:12  */
  assign decimal_exponent = n16537; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:92:12  */
  assign work_mantissa = n16541; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:93:12  */
  assign work_exponent = n16545; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:94:12  */
  assign result_sign = n16549; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:95:12  */
  assign exp_sign = n16553; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:123:12  */
  assign cycle_count = n16555; // (signal)
  /* TG68K_FPU_PackedDecimal.vhd:128:18  */
  always @*
    packed_conversion_temp_mantissa = n16510; // (isignal)
  initial
    packed_conversion_temp_mantissa = 128'bX;
  /* TG68K_FPU_PackedDecimal.vhd:133:19  */
  assign n15692 = ~nreset;
  /* TG68K_FPU_PackedDecimal.vhd:155:25  */
  assign n15695 = start_conversion ? 3'b001 : packed_state;
  /* TG68K_FPU_PackedDecimal.vhd:147:21  */
  assign n15697 = packed_state == 3'b000;
  /* TG68K_FPU_PackedDecimal.vhd:163:53  */
  assign n15698 = packed_in[95]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:164:50  */
  assign n15699 = packed_in[94]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:165:54  */
  assign n15700 = packed_in[91:80]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:166:52  */
  assign n15701 = packed_in[67:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15702 = bcd_digits[3:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15704 = $unsigned(n15702) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15707 = n15704 ? 1'b1 : 1'b0;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15709 = bcd_digits[7:4]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15711 = $unsigned(n15709) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15713 = n15711 ? 1'b1 : n15707;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15714 = bcd_digits[11:8]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15716 = $unsigned(n15714) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15718 = n15716 ? 1'b1 : n15713;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15719 = bcd_digits[15:12]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15721 = $unsigned(n15719) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15723 = n15721 ? 1'b1 : n15718;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15724 = bcd_digits[19:16]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15726 = $unsigned(n15724) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15728 = n15726 ? 1'b1 : n15723;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15729 = bcd_digits[23:20]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15731 = $unsigned(n15729) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15733 = n15731 ? 1'b1 : n15728;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15734 = bcd_digits[27:24]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15736 = $unsigned(n15734) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15738 = n15736 ? 1'b1 : n15733;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15739 = bcd_digits[31:28]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15741 = $unsigned(n15739) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15743 = n15741 ? 1'b1 : n15738;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15744 = bcd_digits[35:32]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15746 = $unsigned(n15744) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15748 = n15746 ? 1'b1 : n15743;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15749 = bcd_digits[39:36]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15751 = $unsigned(n15749) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15753 = n15751 ? 1'b1 : n15748;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15754 = bcd_digits[43:40]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15756 = $unsigned(n15754) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15758 = n15756 ? 1'b1 : n15753;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15759 = bcd_digits[47:44]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15761 = $unsigned(n15759) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15763 = n15761 ? 1'b1 : n15758;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15764 = bcd_digits[51:48]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15766 = $unsigned(n15764) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15768 = n15766 ? 1'b1 : n15763;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15769 = bcd_digits[55:52]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15771 = $unsigned(n15769) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15773 = n15771 ? 1'b1 : n15768;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15774 = bcd_digits[59:56]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15776 = $unsigned(n15774) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15778 = n15776 ? 1'b1 : n15773;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15779 = bcd_digits[63:60]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15781 = $unsigned(n15779) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15783 = n15781 ? 1'b1 : n15778;
  /* TG68K_FPU_PackedDecimal.vhd:171:55  */
  assign n15784 = bcd_digits[67:64]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:171:75  */
  assign n15786 = $unsigned(n15784) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:171:33  */
  assign n15788 = n15786 ? 1'b1 : n15783;
  /* TG68K_FPU_PackedDecimal.vhd:178:57  */
  assign n15789 = bcd_exponent[3:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:178:77  */
  assign n15791 = $unsigned(n15789) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:178:33  */
  assign n15793 = n15791 ? 1'b1 : n15788;
  /* TG68K_FPU_PackedDecimal.vhd:178:57  */
  assign n15794 = bcd_exponent[7:4]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:178:77  */
  assign n15796 = $unsigned(n15794) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:178:33  */
  assign n15798 = n15796 ? 1'b1 : n15793;
  /* TG68K_FPU_PackedDecimal.vhd:178:57  */
  assign n15799 = bcd_exponent[11:8]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:178:77  */
  assign n15801 = $unsigned(n15799) > $unsigned(4'b1001);
  /* TG68K_FPU_PackedDecimal.vhd:178:33  */
  assign n15803 = n15801 ? 1'b1 : n15798;
  /* TG68K_FPU_PackedDecimal.vhd:187:55  */
  assign n15804 = extended_in[79]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:188:77  */
  assign n15805 = extended_in[78:64]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:188:46  */
  assign n15806 = {16'b0, n15805};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:188:94  */
  assign n15807 = {1'b0, n15806};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:188:94  */
  assign n15809 = n15807 - 32'b00000000000000000011111111111111;
  /* TG68K_FPU_PackedDecimal.vhd:189:70  */
  assign n15810 = extended_in[63:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:193:43  */
  assign n15812 = extended_in[78:64]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:193:58  */
  assign n15814 = n15812 == 15'b111111111111111;
  /* TG68K_FPU_PackedDecimal.vhd:195:47  */
  assign n15815 = extended_in[63]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:195:73  */
  assign n15816 = extended_in[62:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:195:87  */
  assign n15818 = n15816 == 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_PackedDecimal.vhd:195:58  */
  assign n15819 = n15818 & n15815;
  /* TG68K_FPU_PackedDecimal.vhd:195:33  */
  assign n15838 = n15819 ? n16563 : 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15840 = n15858 ? 1'b1 : n16565;
  /* TG68K_FPU_PackedDecimal.vhd:195:33  */
  assign n15842 = n15819 ? n16569 : 1'b1;
  /* TG68K_FPU_PackedDecimal.vhd:195:33  */
  assign n15844 = n15819 ? packed_state : 3'b110;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15845 = {4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001};
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15846 = n15861 ? n15845 : bcd_digits;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15848 = n15862 ? 12'b100110011001 : bcd_exponent;
  /* TG68K_FPU_PackedDecimal.vhd:209:46  */
  assign n15849 = extended_in[78:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:209:60  */
  assign n15851 = n15849 == 79'b0000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_PackedDecimal.vhd:209:29  */
  assign n15853 = n15851 ? 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : n16563;
  /* TG68K_FPU_PackedDecimal.vhd:209:29  */
  assign n15856 = n15851 ? 3'b110 : 3'b011;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15857 = n15814 ? n15838 : n15853;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15858 = n15819 & n15814;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15859 = n15814 ? n15842 : n16569;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15860 = n15814 ? n15844 : n15856;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15861 = n15819 & n15814;
  /* TG68K_FPU_PackedDecimal.vhd:193:29  */
  assign n15862 = n15819 & n15814;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15863 = packed_to_extended ? n16563 : n15857;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15864 = packed_to_extended ? n16565 : n15840;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15865 = packed_to_extended ? n15803 : n15859;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15867 = packed_to_extended ? 3'b010 : n15860;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15868 = packed_to_extended ? n15701 : n15846;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15869 = packed_to_extended ? n15700 : n15848;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15870 = {64'b0000000000000000000000000000000000000000000000000000000000000000, n15810};
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15871 = packed_to_extended ? work_mantissa : n15870;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15872 = packed_to_extended ? work_exponent : n15809;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15873 = packed_to_extended ? n15698 : n15804;
  /* TG68K_FPU_PackedDecimal.vhd:160:25  */
  assign n15874 = packed_to_extended ? n15699 : exp_sign;
  /* TG68K_FPU_PackedDecimal.vhd:159:21  */
  assign n15876 = packed_state == 3'b001;
  /* TG68K_FPU_PackedDecimal.vhd:221:40  */
  assign n15877 = {26'b0, cycle_count};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:221:40  */
  assign n15879 = n15877 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_PackedDecimal.vhd:221:25  */
  assign n15881 = n15879 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : binary_mantissa;
  /* TG68K_FPU_PackedDecimal.vhd:221:25  */
  assign n15883 = n15879 ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : packed_conversion_temp_mantissa;
  /* TG68K_FPU_PackedDecimal.vhd:226:40  */
  assign n15884 = {26'b0, cycle_count};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:226:40  */
  assign n15886 = $signed(n15884) < $signed(32'b00000000000000000000000000010001);
  /* TG68K_FPU_PackedDecimal.vhd:229:89  */
  assign n15887 = bcd_digits[67:64]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:229:59  */
  assign n15888 = {27'b0, n15887};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:229:44  */
  assign n15889 = {1'b0, n15888};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:229:33  */
  assign n15891 = cycle_count == 6'b000000;
  /* TG68K_FPU_PackedDecimal.vhd:230:89  */
  assign n15892 = bcd_digits[63:60]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:230:59  */
  assign n15893 = {27'b0, n15892};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:230:44  */
  assign n15894 = {1'b0, n15893};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:230:33  */
  assign n15896 = cycle_count == 6'b000001;
  /* TG68K_FPU_PackedDecimal.vhd:231:89  */
  assign n15897 = bcd_digits[59:56]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:231:59  */
  assign n15898 = {27'b0, n15897};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:231:44  */
  assign n15899 = {1'b0, n15898};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:231:33  */
  assign n15901 = cycle_count == 6'b000010;
  /* TG68K_FPU_PackedDecimal.vhd:232:89  */
  assign n15902 = bcd_digits[55:52]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:232:59  */
  assign n15903 = {27'b0, n15902};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:232:44  */
  assign n15904 = {1'b0, n15903};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:232:33  */
  assign n15906 = cycle_count == 6'b000011;
  /* TG68K_FPU_PackedDecimal.vhd:233:89  */
  assign n15907 = bcd_digits[51:48]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:233:59  */
  assign n15908 = {27'b0, n15907};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:233:44  */
  assign n15909 = {1'b0, n15908};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:233:33  */
  assign n15911 = cycle_count == 6'b000100;
  /* TG68K_FPU_PackedDecimal.vhd:234:89  */
  assign n15912 = bcd_digits[47:44]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:234:59  */
  assign n15913 = {27'b0, n15912};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:234:44  */
  assign n15914 = {1'b0, n15913};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:234:33  */
  assign n15916 = cycle_count == 6'b000101;
  /* TG68K_FPU_PackedDecimal.vhd:235:89  */
  assign n15917 = bcd_digits[43:40]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:235:59  */
  assign n15918 = {27'b0, n15917};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:235:44  */
  assign n15919 = {1'b0, n15918};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:235:33  */
  assign n15921 = cycle_count == 6'b000110;
  /* TG68K_FPU_PackedDecimal.vhd:236:89  */
  assign n15922 = bcd_digits[39:36]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:236:59  */
  assign n15923 = {27'b0, n15922};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:236:44  */
  assign n15924 = {1'b0, n15923};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:236:33  */
  assign n15926 = cycle_count == 6'b000111;
  /* TG68K_FPU_PackedDecimal.vhd:237:89  */
  assign n15927 = bcd_digits[35:32]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:237:59  */
  assign n15928 = {27'b0, n15927};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:237:44  */
  assign n15929 = {1'b0, n15928};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:237:33  */
  assign n15931 = cycle_count == 6'b001000;
  /* TG68K_FPU_PackedDecimal.vhd:238:89  */
  assign n15932 = bcd_digits[31:28]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:238:59  */
  assign n15933 = {27'b0, n15932};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:238:44  */
  assign n15934 = {1'b0, n15933};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:238:33  */
  assign n15936 = cycle_count == 6'b001001;
  /* TG68K_FPU_PackedDecimal.vhd:239:89  */
  assign n15937 = bcd_digits[27:24]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:239:59  */
  assign n15938 = {27'b0, n15937};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:239:44  */
  assign n15939 = {1'b0, n15938};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:239:33  */
  assign n15941 = cycle_count == 6'b001010;
  /* TG68K_FPU_PackedDecimal.vhd:240:89  */
  assign n15942 = bcd_digits[23:20]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:240:59  */
  assign n15943 = {27'b0, n15942};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:240:44  */
  assign n15944 = {1'b0, n15943};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:240:33  */
  assign n15946 = cycle_count == 6'b001011;
  /* TG68K_FPU_PackedDecimal.vhd:241:89  */
  assign n15947 = bcd_digits[19:16]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:241:59  */
  assign n15948 = {27'b0, n15947};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:241:44  */
  assign n15949 = {1'b0, n15948};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:241:33  */
  assign n15951 = cycle_count == 6'b001100;
  /* TG68K_FPU_PackedDecimal.vhd:242:89  */
  assign n15952 = bcd_digits[15:12]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:242:59  */
  assign n15953 = {27'b0, n15952};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:242:44  */
  assign n15954 = {1'b0, n15953};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:242:33  */
  assign n15956 = cycle_count == 6'b001101;
  /* TG68K_FPU_PackedDecimal.vhd:243:89  */
  assign n15957 = bcd_digits[11:8]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:243:59  */
  assign n15958 = {27'b0, n15957};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:243:44  */
  assign n15959 = {1'b0, n15958};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:243:33  */
  assign n15961 = cycle_count == 6'b001110;
  /* TG68K_FPU_PackedDecimal.vhd:244:89  */
  assign n15962 = bcd_digits[7:4]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:244:59  */
  assign n15963 = {27'b0, n15962};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:244:44  */
  assign n15964 = {1'b0, n15963};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:244:33  */
  assign n15966 = cycle_count == 6'b001111;
  /* TG68K_FPU_PackedDecimal.vhd:245:89  */
  assign n15967 = bcd_digits[3:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:245:59  */
  assign n15968 = {27'b0, n15967};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:245:44  */
  assign n15969 = {1'b0, n15968};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:245:33  */
  assign n15971 = cycle_count == 6'b010000;
  /* TG68K_FPU_Exception_Handler.vhd:235:75  */
  assign n15972 = {n15971, n15966, n15961, n15956, n15951, n15946, n15941, n15936, n15931, n15926, n15921, n15916, n15911, n15906, n15901, n15896, n15891};
  /* TG68K_FPU_PackedDecimal.vhd:228:29  */
  always @*
    case (n15972)
      17'b10000000000000000: n15974 = n15969;
      17'b01000000000000000: n15974 = n15964;
      17'b00100000000000000: n15974 = n15959;
      17'b00010000000000000: n15974 = n15954;
      17'b00001000000000000: n15974 = n15949;
      17'b00000100000000000: n15974 = n15944;
      17'b00000010000000000: n15974 = n15939;
      17'b00000001000000000: n15974 = n15934;
      17'b00000000100000000: n15974 = n15929;
      17'b00000000010000000: n15974 = n15924;
      17'b00000000001000000: n15974 = n15919;
      17'b00000000000100000: n15974 = n15914;
      17'b00000000000010000: n15974 = n15909;
      17'b00000000000001000: n15974 = n15904;
      17'b00000000000000100: n15974 = n15899;
      17'b00000000000000010: n15974 = n15894;
      17'b00000000000000001: n15974 = n15889;
      default: n15974 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:249:67  */
  assign n15975 = {128'b0, n15883};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:249:67  */
  assign n15977 = $signed(n15975) * $signed(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010); // smul
  /* TG68K_FPU_PackedDecimal.vhd:249:46  */
  assign n15978 = n15977[127:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:249:78  */
  assign n15979 = n15974[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:249:78  */
  assign n15980 = {97'b0, n15979};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:249:78  */
  assign n15981 = n15978 + n15980;
  /* TG68K_FPU_PackedDecimal.vhd:250:56  */
  assign n15982 = {26'b0, cycle_count};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:250:56  */
  assign n15984 = n15982 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_PackedDecimal.vhd:250:44  */
  assign n15985 = n15984[5:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:101:38  */
  assign n15994 = bcd_exponent[3:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:101:15  */
  assign n15995 = {27'b0, n15994};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:101:9  */
  assign n15996 = {1'b0, n15995};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:102:38  */
  assign n15998 = bcd_exponent[7:4]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:102:15  */
  assign n15999 = {27'b0, n15998};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:102:9  */
  assign n16000 = {1'b0, n15999};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:103:38  */
  assign n16002 = bcd_exponent[11:8]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:103:15  */
  assign n16003 = {27'b0, n16002};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:103:9  */
  assign n16004 = {1'b0, n16003};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:104:15  */
  assign n16007 = $signed(n15996) > $signed(32'b00000000000000000000000000001001);
  /* TG68K_FPU_PackedDecimal.vhd:104:25  */
  assign n16009 = $signed(n16000) > $signed(32'b00000000000000000000000000001001);
  /* TG68K_FPU_PackedDecimal.vhd:104:19  */
  assign n16010 = n16007 | n16009;
  /* TG68K_FPU_PackedDecimal.vhd:104:35  */
  assign n16012 = $signed(n16004) > $signed(32'b00000000000000000000000000001001);
  /* TG68K_FPU_PackedDecimal.vhd:104:29  */
  assign n16013 = n16010 | n16012;
  /* TG68K_FPU_PackedDecimal.vhd:104:9  */
  assign n16017 = n16013 ? 1'b0 : 1'b1;
  /* TG68K_FPU_PackedDecimal.vhd:104:9  */
  assign n16023 = n16013 ? 32'b11111111111111111111111111111111 : 32'bX;
  /* TG68K_FPU_PackedDecimal.vhd:107:19  */
  assign n16025 = $signed(n16004) * $signed(32'b00000000000000000000000001100100); // smul
  /* TG68K_FPU_PackedDecimal.vhd:107:30  */
  assign n16027 = $signed(n16000) * $signed(32'b00000000000000000000000000001010); // smul
  /* TG68K_FPU_PackedDecimal.vhd:107:25  */
  assign n16028 = n16025 + n16027;
  /* TG68K_FPU_PackedDecimal.vhd:107:35  */
  assign n16029 = n16028 + n15996;
  /* TG68K_FPU_PackedDecimal.vhd:107:9  */
  assign n16034 = n16017 ? n16029 : n16023;
  /* TG68K_FPU_PackedDecimal.vhd:254:53  */
  assign n16035 = -n16034;
  /* TG68K_FPU_PackedDecimal.vhd:254:84  */
  assign n16036 = {{25{k_factor[6]}}, k_factor}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:254:82  */
  assign n16037 = n16035 - n16036;
  /* TG68K_FPU_PackedDecimal.vhd:254:53  */
  assign n16038 = n16037[10:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:101:38  */
  assign n16047 = bcd_exponent[3:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:101:15  */
  assign n16048 = {27'b0, n16047};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:101:9  */
  assign n16049 = {1'b0, n16048};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:102:38  */
  assign n16051 = bcd_exponent[7:4]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:102:15  */
  assign n16052 = {27'b0, n16051};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:102:9  */
  assign n16053 = {1'b0, n16052};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:103:38  */
  assign n16055 = bcd_exponent[11:8]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:103:15  */
  assign n16056 = {27'b0, n16055};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:103:9  */
  assign n16057 = {1'b0, n16056};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:104:15  */
  assign n16060 = $signed(n16049) > $signed(32'b00000000000000000000000000001001);
  /* TG68K_FPU_PackedDecimal.vhd:104:25  */
  assign n16062 = $signed(n16053) > $signed(32'b00000000000000000000000000001001);
  /* TG68K_FPU_PackedDecimal.vhd:104:19  */
  assign n16063 = n16060 | n16062;
  /* TG68K_FPU_PackedDecimal.vhd:104:35  */
  assign n16065 = $signed(n16057) > $signed(32'b00000000000000000000000000001001);
  /* TG68K_FPU_PackedDecimal.vhd:104:29  */
  assign n16066 = n16063 | n16065;
  /* TG68K_FPU_PackedDecimal.vhd:104:9  */
  assign n16070 = n16066 ? 1'b0 : 1'b1;
  /* TG68K_FPU_PackedDecimal.vhd:104:9  */
  assign n16076 = n16066 ? 32'b11111111111111111111111111111111 : 32'bX;
  /* TG68K_FPU_PackedDecimal.vhd:107:19  */
  assign n16078 = $signed(n16057) * $signed(32'b00000000000000000000000001100100); // smul
  /* TG68K_FPU_PackedDecimal.vhd:107:30  */
  assign n16080 = $signed(n16053) * $signed(32'b00000000000000000000000000001010); // smul
  /* TG68K_FPU_PackedDecimal.vhd:107:25  */
  assign n16081 = n16078 + n16080;
  /* TG68K_FPU_PackedDecimal.vhd:107:35  */
  assign n16082 = n16081 + n16049;
  /* TG68K_FPU_PackedDecimal.vhd:107:9  */
  assign n16087 = n16070 ? n16082 : n16076;
  /* TG68K_FPU_PackedDecimal.vhd:256:83  */
  assign n16088 = {{25{k_factor[6]}}, k_factor}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:256:81  */
  assign n16089 = n16087 - n16088;
  /* TG68K_FPU_PackedDecimal.vhd:256:53  */
  assign n16090 = n16089[10:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:253:29  */
  assign n16091 = exp_sign ? n16038 : n16090;
  /* TG68K_FPU_PackedDecimal.vhd:259:78  */
  assign n16092 = n15883[63:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:226:25  */
  assign n16094 = n15886 ? packed_state : 3'b100;
  /* TG68K_FPU_PackedDecimal.vhd:226:25  */
  assign n16095 = n15886 ? n15881 : n16092;
  /* TG68K_FPU_PackedDecimal.vhd:226:25  */
  assign n16096 = n15886 ? decimal_exponent : n16091;
  /* TG68K_FPU_PackedDecimal.vhd:226:25  */
  assign n16098 = n15886 ? n15985 : 6'b000000;
  /* TG68K_FPU_PackedDecimal.vhd:226:25  */
  assign n16099 = n15886 ? n15981 : n15883;
  /* TG68K_FPU_PackedDecimal.vhd:218:21  */
  assign n16102 = packed_state == 3'b010;
  /* TG68K_FPU_PackedDecimal.vhd:267:40  */
  assign n16103 = {26'b0, cycle_count};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:267:40  */
  assign n16105 = n16103 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_PackedDecimal.vhd:274:46  */
  assign n16107 = $signed(work_exponent) > $signed(32'b00000000000000000000000000000000);
  /* TG68K_FPU_PackedDecimal.vhd:275:67  */
  assign n16109 = $signed(work_exponent) * $signed(32'b00000000000000000000000000000011); // smul
  /* TG68K_FPU_PackedDecimal.vhd:275:71  */
  assign n16111 = $signed(n16109) / $signed(32'b00000000000000000000000000001010); // sdiv
  /* TG68K_FPU_PackedDecimal.vhd:275:53  */
  assign n16112 = n16111[10:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:278:68  */
  assign n16114 = $signed(work_exponent) * $signed(32'b00000000000000000000000000000011); // smul
  /* TG68K_FPU_PackedDecimal.vhd:278:72  */
  assign n16116 = $signed(n16114) / $signed(32'b00000000000000000000000000001010); // sdiv
  /* TG68K_FPU_PackedDecimal.vhd:278:53  */
  assign n16117 = -n16116;
  /* TG68K_FPU_PackedDecimal.vhd:278:53  */
  assign n16118 = n16117[10:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:274:29  */
  assign n16119 = n16107 ? n16112 : n16118;
  /* TG68K_FPU_PackedDecimal.vhd:274:29  */
  assign n16122 = n16107 ? 1'b0 : 1'b1;
  /* TG68K_FPU_PackedDecimal.vhd:267:25  */
  assign n16124 = n16105 ? 68'b00000000000000000000000000000000000000000000000000000000000000000000 : bcd_digits;
  /* TG68K_FPU_PackedDecimal.vhd:267:25  */
  assign n16125 = n16105 ? n16119 : decimal_exponent;
  /* TG68K_FPU_PackedDecimal.vhd:267:25  */
  assign n16126 = n16105 ? n16122 : exp_sign;
  /* TG68K_FPU_PackedDecimal.vhd:267:25  */
  assign n16127 = n16105 ? work_mantissa : packed_conversion_temp_mantissa;
  /* TG68K_FPU_PackedDecimal.vhd:283:40  */
  assign n16128 = {26'b0, cycle_count};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:283:40  */
  assign n16130 = $signed(n16128) < $signed(32'b00000000000000000000000000010001);
  /* TG68K_FPU_PackedDecimal.vhd:286:102  */
  assign n16131 = n16127[3:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:286:115  */
  assign n16133 = n16131 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:286:33  */
  assign n16135 = cycle_count == 6'b000000;
  /* TG68K_FPU_PackedDecimal.vhd:287:102  */
  assign n16136 = n16127[7:4]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:287:115  */
  assign n16138 = n16136 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:287:33  */
  assign n16140 = cycle_count == 6'b000001;
  /* TG68K_FPU_PackedDecimal.vhd:288:102  */
  assign n16141 = n16127[11:8]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:288:116  */
  assign n16143 = n16141 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:288:33  */
  assign n16145 = cycle_count == 6'b000010;
  /* TG68K_FPU_PackedDecimal.vhd:289:102  */
  assign n16146 = n16127[15:12]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:289:117  */
  assign n16148 = n16146 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:289:33  */
  assign n16150 = cycle_count == 6'b000011;
  /* TG68K_FPU_PackedDecimal.vhd:290:102  */
  assign n16151 = n16127[19:16]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:290:117  */
  assign n16153 = n16151 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:290:33  */
  assign n16155 = cycle_count == 6'b000100;
  /* TG68K_FPU_PackedDecimal.vhd:291:102  */
  assign n16156 = n16127[23:20]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:291:117  */
  assign n16158 = n16156 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:291:33  */
  assign n16160 = cycle_count == 6'b000101;
  /* TG68K_FPU_PackedDecimal.vhd:292:102  */
  assign n16161 = n16127[27:24]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:292:117  */
  assign n16163 = n16161 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:292:33  */
  assign n16165 = cycle_count == 6'b000110;
  /* TG68K_FPU_PackedDecimal.vhd:293:102  */
  assign n16166 = n16127[31:28]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:293:117  */
  assign n16168 = n16166 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:293:33  */
  assign n16170 = cycle_count == 6'b000111;
  /* TG68K_FPU_PackedDecimal.vhd:294:102  */
  assign n16171 = n16127[35:32]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:294:117  */
  assign n16173 = n16171 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:294:33  */
  assign n16175 = cycle_count == 6'b001000;
  /* TG68K_FPU_PackedDecimal.vhd:295:102  */
  assign n16176 = n16127[39:36]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:295:117  */
  assign n16178 = n16176 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:295:33  */
  assign n16180 = cycle_count == 6'b001001;
  /* TG68K_FPU_PackedDecimal.vhd:296:102  */
  assign n16181 = n16127[43:40]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:296:117  */
  assign n16183 = n16181 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:296:33  */
  assign n16185 = cycle_count == 6'b001010;
  /* TG68K_FPU_PackedDecimal.vhd:297:102  */
  assign n16186 = n16127[47:44]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:297:117  */
  assign n16188 = n16186 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:297:33  */
  assign n16190 = cycle_count == 6'b001011;
  /* TG68K_FPU_PackedDecimal.vhd:298:102  */
  assign n16191 = n16127[51:48]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:298:117  */
  assign n16193 = n16191 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:298:33  */
  assign n16195 = cycle_count == 6'b001100;
  /* TG68K_FPU_PackedDecimal.vhd:299:102  */
  assign n16196 = n16127[55:52]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:299:117  */
  assign n16198 = n16196 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:299:33  */
  assign n16200 = cycle_count == 6'b001101;
  /* TG68K_FPU_PackedDecimal.vhd:300:102  */
  assign n16201 = n16127[59:56]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:300:117  */
  assign n16203 = n16201 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:300:33  */
  assign n16205 = cycle_count == 6'b001110;
  /* TG68K_FPU_PackedDecimal.vhd:301:102  */
  assign n16206 = n16127[63:60]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:301:117  */
  assign n16208 = n16206 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:301:33  */
  assign n16210 = cycle_count == 6'b001111;
  /* TG68K_FPU_PackedDecimal.vhd:302:102  */
  assign n16211 = n16127[67:64]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:302:117  */
  assign n16213 = n16211 & 4'b1001;
  /* TG68K_FPU_PackedDecimal.vhd:302:33  */
  assign n16215 = cycle_count == 6'b010000;
  assign n16216 = {n16215, n16210, n16205, n16200, n16195, n16190, n16185, n16180, n16175, n16170, n16165, n16160, n16155, n16150, n16145, n16140, n16135};
  assign n16217 = n16124[3:0]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16218 = n16217;
      17'b01000000000000000: n16218 = n16217;
      17'b00100000000000000: n16218 = n16217;
      17'b00010000000000000: n16218 = n16217;
      17'b00001000000000000: n16218 = n16217;
      17'b00000100000000000: n16218 = n16217;
      17'b00000010000000000: n16218 = n16217;
      17'b00000001000000000: n16218 = n16217;
      17'b00000000100000000: n16218 = n16217;
      17'b00000000010000000: n16218 = n16217;
      17'b00000000001000000: n16218 = n16217;
      17'b00000000000100000: n16218 = n16217;
      17'b00000000000010000: n16218 = n16217;
      17'b00000000000001000: n16218 = n16217;
      17'b00000000000000100: n16218 = n16217;
      17'b00000000000000010: n16218 = n16217;
      17'b00000000000000001: n16218 = n16133;
      default: n16218 = n16217;
    endcase
  assign n16219 = n16124[7:4]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16220 = n16219;
      17'b01000000000000000: n16220 = n16219;
      17'b00100000000000000: n16220 = n16219;
      17'b00010000000000000: n16220 = n16219;
      17'b00001000000000000: n16220 = n16219;
      17'b00000100000000000: n16220 = n16219;
      17'b00000010000000000: n16220 = n16219;
      17'b00000001000000000: n16220 = n16219;
      17'b00000000100000000: n16220 = n16219;
      17'b00000000010000000: n16220 = n16219;
      17'b00000000001000000: n16220 = n16219;
      17'b00000000000100000: n16220 = n16219;
      17'b00000000000010000: n16220 = n16219;
      17'b00000000000001000: n16220 = n16219;
      17'b00000000000000100: n16220 = n16219;
      17'b00000000000000010: n16220 = n16138;
      17'b00000000000000001: n16220 = n16219;
      default: n16220 = n16219;
    endcase
  assign n16221 = n16124[11:8]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16222 = n16221;
      17'b01000000000000000: n16222 = n16221;
      17'b00100000000000000: n16222 = n16221;
      17'b00010000000000000: n16222 = n16221;
      17'b00001000000000000: n16222 = n16221;
      17'b00000100000000000: n16222 = n16221;
      17'b00000010000000000: n16222 = n16221;
      17'b00000001000000000: n16222 = n16221;
      17'b00000000100000000: n16222 = n16221;
      17'b00000000010000000: n16222 = n16221;
      17'b00000000001000000: n16222 = n16221;
      17'b00000000000100000: n16222 = n16221;
      17'b00000000000010000: n16222 = n16221;
      17'b00000000000001000: n16222 = n16221;
      17'b00000000000000100: n16222 = n16143;
      17'b00000000000000010: n16222 = n16221;
      17'b00000000000000001: n16222 = n16221;
      default: n16222 = n16221;
    endcase
  assign n16223 = n16124[15:12]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16224 = n16223;
      17'b01000000000000000: n16224 = n16223;
      17'b00100000000000000: n16224 = n16223;
      17'b00010000000000000: n16224 = n16223;
      17'b00001000000000000: n16224 = n16223;
      17'b00000100000000000: n16224 = n16223;
      17'b00000010000000000: n16224 = n16223;
      17'b00000001000000000: n16224 = n16223;
      17'b00000000100000000: n16224 = n16223;
      17'b00000000010000000: n16224 = n16223;
      17'b00000000001000000: n16224 = n16223;
      17'b00000000000100000: n16224 = n16223;
      17'b00000000000010000: n16224 = n16223;
      17'b00000000000001000: n16224 = n16148;
      17'b00000000000000100: n16224 = n16223;
      17'b00000000000000010: n16224 = n16223;
      17'b00000000000000001: n16224 = n16223;
      default: n16224 = n16223;
    endcase
  assign n16225 = n16124[19:16]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16226 = n16225;
      17'b01000000000000000: n16226 = n16225;
      17'b00100000000000000: n16226 = n16225;
      17'b00010000000000000: n16226 = n16225;
      17'b00001000000000000: n16226 = n16225;
      17'b00000100000000000: n16226 = n16225;
      17'b00000010000000000: n16226 = n16225;
      17'b00000001000000000: n16226 = n16225;
      17'b00000000100000000: n16226 = n16225;
      17'b00000000010000000: n16226 = n16225;
      17'b00000000001000000: n16226 = n16225;
      17'b00000000000100000: n16226 = n16225;
      17'b00000000000010000: n16226 = n16153;
      17'b00000000000001000: n16226 = n16225;
      17'b00000000000000100: n16226 = n16225;
      17'b00000000000000010: n16226 = n16225;
      17'b00000000000000001: n16226 = n16225;
      default: n16226 = n16225;
    endcase
  assign n16227 = n16124[23:20]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16228 = n16227;
      17'b01000000000000000: n16228 = n16227;
      17'b00100000000000000: n16228 = n16227;
      17'b00010000000000000: n16228 = n16227;
      17'b00001000000000000: n16228 = n16227;
      17'b00000100000000000: n16228 = n16227;
      17'b00000010000000000: n16228 = n16227;
      17'b00000001000000000: n16228 = n16227;
      17'b00000000100000000: n16228 = n16227;
      17'b00000000010000000: n16228 = n16227;
      17'b00000000001000000: n16228 = n16227;
      17'b00000000000100000: n16228 = n16158;
      17'b00000000000010000: n16228 = n16227;
      17'b00000000000001000: n16228 = n16227;
      17'b00000000000000100: n16228 = n16227;
      17'b00000000000000010: n16228 = n16227;
      17'b00000000000000001: n16228 = n16227;
      default: n16228 = n16227;
    endcase
  assign n16229 = n16124[27:24]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16230 = n16229;
      17'b01000000000000000: n16230 = n16229;
      17'b00100000000000000: n16230 = n16229;
      17'b00010000000000000: n16230 = n16229;
      17'b00001000000000000: n16230 = n16229;
      17'b00000100000000000: n16230 = n16229;
      17'b00000010000000000: n16230 = n16229;
      17'b00000001000000000: n16230 = n16229;
      17'b00000000100000000: n16230 = n16229;
      17'b00000000010000000: n16230 = n16229;
      17'b00000000001000000: n16230 = n16163;
      17'b00000000000100000: n16230 = n16229;
      17'b00000000000010000: n16230 = n16229;
      17'b00000000000001000: n16230 = n16229;
      17'b00000000000000100: n16230 = n16229;
      17'b00000000000000010: n16230 = n16229;
      17'b00000000000000001: n16230 = n16229;
      default: n16230 = n16229;
    endcase
  assign n16231 = n16124[31:28]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16232 = n16231;
      17'b01000000000000000: n16232 = n16231;
      17'b00100000000000000: n16232 = n16231;
      17'b00010000000000000: n16232 = n16231;
      17'b00001000000000000: n16232 = n16231;
      17'b00000100000000000: n16232 = n16231;
      17'b00000010000000000: n16232 = n16231;
      17'b00000001000000000: n16232 = n16231;
      17'b00000000100000000: n16232 = n16231;
      17'b00000000010000000: n16232 = n16168;
      17'b00000000001000000: n16232 = n16231;
      17'b00000000000100000: n16232 = n16231;
      17'b00000000000010000: n16232 = n16231;
      17'b00000000000001000: n16232 = n16231;
      17'b00000000000000100: n16232 = n16231;
      17'b00000000000000010: n16232 = n16231;
      17'b00000000000000001: n16232 = n16231;
      default: n16232 = n16231;
    endcase
  assign n16233 = n16124[35:32]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16234 = n16233;
      17'b01000000000000000: n16234 = n16233;
      17'b00100000000000000: n16234 = n16233;
      17'b00010000000000000: n16234 = n16233;
      17'b00001000000000000: n16234 = n16233;
      17'b00000100000000000: n16234 = n16233;
      17'b00000010000000000: n16234 = n16233;
      17'b00000001000000000: n16234 = n16233;
      17'b00000000100000000: n16234 = n16173;
      17'b00000000010000000: n16234 = n16233;
      17'b00000000001000000: n16234 = n16233;
      17'b00000000000100000: n16234 = n16233;
      17'b00000000000010000: n16234 = n16233;
      17'b00000000000001000: n16234 = n16233;
      17'b00000000000000100: n16234 = n16233;
      17'b00000000000000010: n16234 = n16233;
      17'b00000000000000001: n16234 = n16233;
      default: n16234 = n16233;
    endcase
  assign n16235 = n16124[39:36]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16236 = n16235;
      17'b01000000000000000: n16236 = n16235;
      17'b00100000000000000: n16236 = n16235;
      17'b00010000000000000: n16236 = n16235;
      17'b00001000000000000: n16236 = n16235;
      17'b00000100000000000: n16236 = n16235;
      17'b00000010000000000: n16236 = n16235;
      17'b00000001000000000: n16236 = n16178;
      17'b00000000100000000: n16236 = n16235;
      17'b00000000010000000: n16236 = n16235;
      17'b00000000001000000: n16236 = n16235;
      17'b00000000000100000: n16236 = n16235;
      17'b00000000000010000: n16236 = n16235;
      17'b00000000000001000: n16236 = n16235;
      17'b00000000000000100: n16236 = n16235;
      17'b00000000000000010: n16236 = n16235;
      17'b00000000000000001: n16236 = n16235;
      default: n16236 = n16235;
    endcase
  assign n16237 = n16124[43:40]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16238 = n16237;
      17'b01000000000000000: n16238 = n16237;
      17'b00100000000000000: n16238 = n16237;
      17'b00010000000000000: n16238 = n16237;
      17'b00001000000000000: n16238 = n16237;
      17'b00000100000000000: n16238 = n16237;
      17'b00000010000000000: n16238 = n16183;
      17'b00000001000000000: n16238 = n16237;
      17'b00000000100000000: n16238 = n16237;
      17'b00000000010000000: n16238 = n16237;
      17'b00000000001000000: n16238 = n16237;
      17'b00000000000100000: n16238 = n16237;
      17'b00000000000010000: n16238 = n16237;
      17'b00000000000001000: n16238 = n16237;
      17'b00000000000000100: n16238 = n16237;
      17'b00000000000000010: n16238 = n16237;
      17'b00000000000000001: n16238 = n16237;
      default: n16238 = n16237;
    endcase
  assign n16239 = n16124[47:44]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16240 = n16239;
      17'b01000000000000000: n16240 = n16239;
      17'b00100000000000000: n16240 = n16239;
      17'b00010000000000000: n16240 = n16239;
      17'b00001000000000000: n16240 = n16239;
      17'b00000100000000000: n16240 = n16188;
      17'b00000010000000000: n16240 = n16239;
      17'b00000001000000000: n16240 = n16239;
      17'b00000000100000000: n16240 = n16239;
      17'b00000000010000000: n16240 = n16239;
      17'b00000000001000000: n16240 = n16239;
      17'b00000000000100000: n16240 = n16239;
      17'b00000000000010000: n16240 = n16239;
      17'b00000000000001000: n16240 = n16239;
      17'b00000000000000100: n16240 = n16239;
      17'b00000000000000010: n16240 = n16239;
      17'b00000000000000001: n16240 = n16239;
      default: n16240 = n16239;
    endcase
  assign n16241 = n16124[51:48]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16242 = n16241;
      17'b01000000000000000: n16242 = n16241;
      17'b00100000000000000: n16242 = n16241;
      17'b00010000000000000: n16242 = n16241;
      17'b00001000000000000: n16242 = n16193;
      17'b00000100000000000: n16242 = n16241;
      17'b00000010000000000: n16242 = n16241;
      17'b00000001000000000: n16242 = n16241;
      17'b00000000100000000: n16242 = n16241;
      17'b00000000010000000: n16242 = n16241;
      17'b00000000001000000: n16242 = n16241;
      17'b00000000000100000: n16242 = n16241;
      17'b00000000000010000: n16242 = n16241;
      17'b00000000000001000: n16242 = n16241;
      17'b00000000000000100: n16242 = n16241;
      17'b00000000000000010: n16242 = n16241;
      17'b00000000000000001: n16242 = n16241;
      default: n16242 = n16241;
    endcase
  assign n16243 = n16124[55:52]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16244 = n16243;
      17'b01000000000000000: n16244 = n16243;
      17'b00100000000000000: n16244 = n16243;
      17'b00010000000000000: n16244 = n16198;
      17'b00001000000000000: n16244 = n16243;
      17'b00000100000000000: n16244 = n16243;
      17'b00000010000000000: n16244 = n16243;
      17'b00000001000000000: n16244 = n16243;
      17'b00000000100000000: n16244 = n16243;
      17'b00000000010000000: n16244 = n16243;
      17'b00000000001000000: n16244 = n16243;
      17'b00000000000100000: n16244 = n16243;
      17'b00000000000010000: n16244 = n16243;
      17'b00000000000001000: n16244 = n16243;
      17'b00000000000000100: n16244 = n16243;
      17'b00000000000000010: n16244 = n16243;
      17'b00000000000000001: n16244 = n16243;
      default: n16244 = n16243;
    endcase
  assign n16245 = n16124[59:56]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16246 = n16245;
      17'b01000000000000000: n16246 = n16245;
      17'b00100000000000000: n16246 = n16203;
      17'b00010000000000000: n16246 = n16245;
      17'b00001000000000000: n16246 = n16245;
      17'b00000100000000000: n16246 = n16245;
      17'b00000010000000000: n16246 = n16245;
      17'b00000001000000000: n16246 = n16245;
      17'b00000000100000000: n16246 = n16245;
      17'b00000000010000000: n16246 = n16245;
      17'b00000000001000000: n16246 = n16245;
      17'b00000000000100000: n16246 = n16245;
      17'b00000000000010000: n16246 = n16245;
      17'b00000000000001000: n16246 = n16245;
      17'b00000000000000100: n16246 = n16245;
      17'b00000000000000010: n16246 = n16245;
      17'b00000000000000001: n16246 = n16245;
      default: n16246 = n16245;
    endcase
  assign n16247 = n16124[63:60]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16248 = n16247;
      17'b01000000000000000: n16248 = n16208;
      17'b00100000000000000: n16248 = n16247;
      17'b00010000000000000: n16248 = n16247;
      17'b00001000000000000: n16248 = n16247;
      17'b00000100000000000: n16248 = n16247;
      17'b00000010000000000: n16248 = n16247;
      17'b00000001000000000: n16248 = n16247;
      17'b00000000100000000: n16248 = n16247;
      17'b00000000010000000: n16248 = n16247;
      17'b00000000001000000: n16248 = n16247;
      17'b00000000000100000: n16248 = n16247;
      17'b00000000000010000: n16248 = n16247;
      17'b00000000000001000: n16248 = n16247;
      17'b00000000000000100: n16248 = n16247;
      17'b00000000000000010: n16248 = n16247;
      17'b00000000000000001: n16248 = n16247;
      default: n16248 = n16247;
    endcase
  assign n16249 = n16124[67:64]; // extract
  /* TG68K_FPU_PackedDecimal.vhd:285:29  */
  always @*
    case (n16216)
      17'b10000000000000000: n16250 = n16213;
      17'b01000000000000000: n16250 = n16249;
      17'b00100000000000000: n16250 = n16249;
      17'b00010000000000000: n16250 = n16249;
      17'b00001000000000000: n16250 = n16249;
      17'b00000100000000000: n16250 = n16249;
      17'b00000010000000000: n16250 = n16249;
      17'b00000001000000000: n16250 = n16249;
      17'b00000000100000000: n16250 = n16249;
      17'b00000000010000000: n16250 = n16249;
      17'b00000000001000000: n16250 = n16249;
      17'b00000000000100000: n16250 = n16249;
      17'b00000000000010000: n16250 = n16249;
      17'b00000000000001000: n16250 = n16249;
      17'b00000000000000100: n16250 = n16249;
      17'b00000000000000010: n16250 = n16249;
      17'b00000000000000001: n16250 = n16249;
      default: n16250 = n16249;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:305:56  */
  assign n16251 = {26'b0, cycle_count};  //  uext
  /* TG68K_FPU_PackedDecimal.vhd:305:56  */
  assign n16253 = n16251 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_PackedDecimal.vhd:305:44  */
  assign n16254 = n16253[5:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:308:66  */
  assign n16255 = {{21{decimal_exponent[10]}}, decimal_exponent}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:308:68  */
  assign n16256 = {{25{k_factor[6]}}, k_factor}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:308:66  */
  assign n16257 = n16255 + n16256;
  /* TG68K_FPU_PackedDecimal.vhd:308:49  */
  assign n16258 = n16257[10:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:311:49  */
  assign n16259 = {{21{decimal_exponent[10]}}, decimal_exponent}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:311:49  */
  assign n16261 = $signed(n16259) < $signed(32'b00000000000000000000000000000000);
  /* TG68K_FPU_PackedDecimal.vhd:313:63  */
  assign n16263 = {{21{decimal_exponent[10]}}, decimal_exponent}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:313:63  */
  assign n16264 = -n16263;
  /* TG68K_FPU_PackedDecimal.vhd:114:65  */
  assign n16271 = n16264 % 32'b00000000000000000000000000001010; // smod
  /* TG68K_FPU_PackedDecimal.vhd:114:60  */
  assign n16272 = n16271[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:114:48  */
  assign n16273 = n16272[3:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:115:22  */
  assign n16277 = $signed(n16264) / $signed(32'b00000000000000000000000000001010); // sdiv
  /* TG68K_FPU_PackedDecimal.vhd:116:65  */
  assign n16279 = n16277 % 32'b00000000000000000000000000001010; // smod
  /* TG68K_FPU_PackedDecimal.vhd:116:60  */
  assign n16280 = n16279[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:116:48  */
  assign n16281 = n16280[3:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:117:22  */
  assign n16284 = $signed(n16277) / $signed(32'b00000000000000000000000000001010); // sdiv
  /* TG68K_FPU_PackedDecimal.vhd:118:66  */
  assign n16286 = n16284 % 32'b00000000000000000000000000001010; // smod
  /* TG68K_FPU_PackedDecimal.vhd:118:61  */
  assign n16287 = n16286[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:118:49  */
  assign n16288 = n16287[3:0];  // trunc
  assign n16289 = {n16288, n16281, n16273};
  /* TG68K_FPU_PackedDecimal.vhd:316:63  */
  assign n16291 = {{21{decimal_exponent[10]}}, decimal_exponent}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:114:65  */
  assign n16298 = n16291 % 32'b00000000000000000000000000001010; // smod
  /* TG68K_FPU_PackedDecimal.vhd:114:60  */
  assign n16299 = n16298[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:114:48  */
  assign n16300 = n16299[3:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:115:22  */
  assign n16304 = $signed(n16291) / $signed(32'b00000000000000000000000000001010); // sdiv
  /* TG68K_FPU_PackedDecimal.vhd:116:65  */
  assign n16306 = n16304 % 32'b00000000000000000000000000001010; // smod
  /* TG68K_FPU_PackedDecimal.vhd:116:60  */
  assign n16307 = n16306[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:116:48  */
  assign n16308 = n16307[3:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:117:22  */
  assign n16311 = $signed(n16304) / $signed(32'b00000000000000000000000000001010); // sdiv
  /* TG68K_FPU_PackedDecimal.vhd:118:66  */
  assign n16313 = n16311 % 32'b00000000000000000000000000001010; // smod
  /* TG68K_FPU_PackedDecimal.vhd:118:61  */
  assign n16314 = n16313[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:118:49  */
  assign n16315 = n16314[3:0];  // trunc
  assign n16316 = {n16315, n16308, n16300};
  /* TG68K_FPU_PackedDecimal.vhd:311:29  */
  assign n16317 = n16261 ? n16289 : n16316;
  /* TG68K_FPU_PackedDecimal.vhd:311:29  */
  assign n16320 = n16261 ? 1'b1 : 1'b0;
  /* TG68K_FPU_PackedDecimal.vhd:283:25  */
  assign n16322 = n16130 ? n16567 : 1'b1;
  /* TG68K_FPU_PackedDecimal.vhd:283:25  */
  assign n16324 = n16130 ? packed_state : 3'b110;
  assign n16325 = {n16250, n16248, n16246, n16244, n16242, n16240, n16238, n16236, n16234, n16232, n16230, n16228, n16226, n16224, n16222, n16220, n16218};
  /* TG68K_FPU_PackedDecimal.vhd:283:25  */
  assign n16326 = n16130 ? n16325 : n16124;
  /* TG68K_FPU_PackedDecimal.vhd:283:25  */
  assign n16327 = n16130 ? bcd_exponent : n16317;
  /* TG68K_FPU_PackedDecimal.vhd:283:25  */
  assign n16328 = n16130 ? n16125 : n16258;
  /* TG68K_FPU_PackedDecimal.vhd:283:25  */
  assign n16329 = n16130 ? n16126 : n16320;
  /* TG68K_FPU_PackedDecimal.vhd:283:25  */
  assign n16330 = n16130 ? n16254 : cycle_count;
  /* TG68K_FPU_PackedDecimal.vhd:264:21  */
  assign n16332 = packed_state == 3'b011;
  /* TG68K_FPU_PackedDecimal.vhd:325:44  */
  assign n16334 = binary_mantissa == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_PackedDecimal.vhd:331:58  */
  assign n16335 = {{21{decimal_exponent[10]}}, decimal_exponent}; // sext
  /* TG68K_FPU_PackedDecimal.vhd:331:58  */
  assign n16337 = $signed(n16335) * $signed(32'b00000000000000000000000000001010); // smul
  /* TG68K_FPU_PackedDecimal.vhd:331:63  */
  assign n16339 = $signed(n16337) / $signed(32'b00000000000000000000000000000011); // sdiv
  /* TG68K_FPU_PackedDecimal.vhd:331:67  */
  assign n16341 = n16339 + 32'b00000000000000000011111111111111;
  /* TG68K_FPU_PackedDecimal.vhd:333:41  */
  assign n16343 = $signed(n16341) < $signed(32'b00000000000000000000000000000000);
  /* TG68K_FPU_PackedDecimal.vhd:335:61  */
  assign n16345 = {result_sign, 79'b0000000000000000000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU_PackedDecimal.vhd:336:44  */
  assign n16347 = $signed(n16341) > $signed(32'b00000000000000000111111111111111);
  /* TG68K_FPU_PackedDecimal.vhd:339:61  */
  assign n16349 = {result_sign, 15'b111111111111111};
  /* TG68K_FPU_PackedDecimal.vhd:339:81  */
  assign n16351 = {n16349, 1'b1};
  /* TG68K_FPU_PackedDecimal.vhd:339:87  */
  assign n16353 = {n16351, 63'b000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU_PackedDecimal.vhd:342:92  */
  assign n16354 = n16341[30:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:342:80  */
  assign n16355 = n16354[14:0];  // trunc
  /* TG68K_FPU_PackedDecimal.vhd:342:61  */
  assign n16356 = {result_sign, n16355};
  /* TG68K_FPU_PackedDecimal.vhd:342:107  */
  assign n16357 = {n16356, binary_mantissa};
  /* TG68K_FPU_PackedDecimal.vhd:336:29  */
  assign n16358 = n16347 ? n16353 : n16357;
  /* TG68K_FPU_PackedDecimal.vhd:336:29  */
  assign n16360 = n16347 ? 1'b1 : n16565;
  /* TG68K_FPU_PackedDecimal.vhd:333:29  */
  assign n16361 = n16343 ? n16345 : n16358;
  /* TG68K_FPU_PackedDecimal.vhd:333:29  */
  assign n16362 = n16343 ? n16565 : n16360;
  /* TG68K_FPU_PackedDecimal.vhd:325:25  */
  assign n16364 = n16334 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n16361;
  /* TG68K_FPU_PackedDecimal.vhd:325:25  */
  assign n16365 = n16334 ? n16565 : n16362;
  /* TG68K_FPU_PackedDecimal.vhd:323:21  */
  assign n16368 = packed_state == 3'b100;
  /* TG68K_FPU_PackedDecimal.vhd:348:21  */
  assign n16370 = packed_state == 3'b101;
  /* TG68K_FPU_PackedDecimal.vhd:354:47  */
  assign n16371 = ~packed_to_extended;
  /* TG68K_FPU_PackedDecimal.vhd:356:55  */
  assign n16372 = {result_sign, exp_sign};
  /* TG68K_FPU_PackedDecimal.vhd:356:66  */
  assign n16374 = {n16372, 2'b00};
  /* TG68K_FPU_PackedDecimal.vhd:356:73  */
  assign n16375 = {n16374, bcd_exponent};
  /* TG68K_FPU_PackedDecimal.vhd:356:88  */
  assign n16377 = {n16375, 1'b0};
  /* TG68K_FPU_PackedDecimal.vhd:356:94  */
  assign n16379 = {n16377, 11'b00000000000};
  /* TG68K_FPU_PackedDecimal.vhd:356:110  */
  assign n16380 = {n16379, bcd_digits};
  /* TG68K_FPU_PackedDecimal.vhd:354:25  */
  assign n16381 = n16371 ? n16380 : n16563;
  /* TG68K_FPU_PackedDecimal.vhd:353:21  */
  assign n16383 = packed_state == 3'b110;
  assign n16384 = {n16383, n16370, n16368, n16332, n16102, n15876, n15697};
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16388 = 1'b1;
      7'b0100000: n16388 = n16557;
      7'b0010000: n16388 = n16557;
      7'b0001000: n16388 = n16557;
      7'b0000100: n16388 = n16557;
      7'b0000010: n16388 = n16557;
      7'b0000001: n16388 = 1'b0;
      default: n16388 = 1'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16392 = 1'b1;
      7'b0100000: n16392 = n16559;
      7'b0010000: n16392 = n16559;
      7'b0001000: n16392 = n16559;
      7'b0000100: n16392 = n16559;
      7'b0000010: n16392 = n16559;
      7'b0000001: n16392 = 1'b0;
      default: n16392 = 1'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16394 = n16561;
      7'b0100000: n16394 = n16561;
      7'b0010000: n16394 = n16364;
      7'b0001000: n16394 = n16561;
      7'b0000100: n16394 = n16561;
      7'b0000010: n16394 = n16561;
      7'b0000001: n16394 = n16561;
      default: n16394 = 80'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16396 = n16381;
      7'b0100000: n16396 = n16563;
      7'b0010000: n16396 = n16563;
      7'b0001000: n16396 = n16563;
      7'b0000100: n16396 = n16563;
      7'b0000010: n16396 = n15863;
      7'b0000001: n16396 = n16563;
      default: n16396 = 96'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16399 = n16565;
      7'b0100000: n16399 = n16565;
      7'b0010000: n16399 = n16365;
      7'b0001000: n16399 = n16565;
      7'b0000100: n16399 = n16565;
      7'b0000010: n16399 = n15864;
      7'b0000001: n16399 = 1'b0;
      default: n16399 = 1'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16403 = n16567;
      7'b0100000: n16403 = n16567;
      7'b0010000: n16403 = 1'b1;
      7'b0001000: n16403 = n16322;
      7'b0000100: n16403 = n16567;
      7'b0000010: n16403 = n16567;
      7'b0000001: n16403 = 1'b0;
      default: n16403 = 1'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16406 = n16569;
      7'b0100000: n16406 = n16569;
      7'b0010000: n16406 = n16569;
      7'b0001000: n16406 = n16569;
      7'b0000100: n16406 = n16569;
      7'b0000010: n16406 = n15865;
      7'b0000001: n16406 = 1'b0;
      default: n16406 = 1'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16411 = 3'b000;
      7'b0100000: n16411 = 3'b110;
      7'b0010000: n16411 = 3'b110;
      7'b0001000: n16411 = n16324;
      7'b0000100: n16411 = n16094;
      7'b0000010: n16411 = n15867;
      7'b0000001: n16411 = n15695;
      default: n16411 = 3'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16413 = bcd_digits;
      7'b0100000: n16413 = bcd_digits;
      7'b0010000: n16413 = bcd_digits;
      7'b0001000: n16413 = n16326;
      7'b0000100: n16413 = bcd_digits;
      7'b0000010: n16413 = n15868;
      7'b0000001: n16413 = bcd_digits;
      default: n16413 = 68'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16415 = bcd_exponent;
      7'b0100000: n16415 = bcd_exponent;
      7'b0010000: n16415 = bcd_exponent;
      7'b0001000: n16415 = n16327;
      7'b0000100: n16415 = bcd_exponent;
      7'b0000010: n16415 = n15869;
      7'b0000001: n16415 = bcd_exponent;
      default: n16415 = 12'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16417 = binary_mantissa;
      7'b0100000: n16417 = binary_mantissa;
      7'b0010000: n16417 = binary_mantissa;
      7'b0001000: n16417 = binary_mantissa;
      7'b0000100: n16417 = n16095;
      7'b0000010: n16417 = binary_mantissa;
      7'b0000001: n16417 = binary_mantissa;
      default: n16417 = 64'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16419 = decimal_exponent;
      7'b0100000: n16419 = decimal_exponent;
      7'b0010000: n16419 = decimal_exponent;
      7'b0001000: n16419 = n16328;
      7'b0000100: n16419 = n16096;
      7'b0000010: n16419 = decimal_exponent;
      7'b0000001: n16419 = decimal_exponent;
      default: n16419 = 11'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16421 = work_mantissa;
      7'b0100000: n16421 = work_mantissa;
      7'b0010000: n16421 = work_mantissa;
      7'b0001000: n16421 = work_mantissa;
      7'b0000100: n16421 = work_mantissa;
      7'b0000010: n16421 = n15871;
      7'b0000001: n16421 = work_mantissa;
      default: n16421 = 128'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16423 = work_exponent;
      7'b0100000: n16423 = work_exponent;
      7'b0010000: n16423 = work_exponent;
      7'b0001000: n16423 = work_exponent;
      7'b0000100: n16423 = work_exponent;
      7'b0000010: n16423 = n15872;
      7'b0000001: n16423 = work_exponent;
      default: n16423 = 32'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16425 = result_sign;
      7'b0100000: n16425 = result_sign;
      7'b0010000: n16425 = result_sign;
      7'b0001000: n16425 = result_sign;
      7'b0000100: n16425 = result_sign;
      7'b0000010: n16425 = n15873;
      7'b0000001: n16425 = result_sign;
      default: n16425 = 1'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16427 = exp_sign;
      7'b0100000: n16427 = exp_sign;
      7'b0010000: n16427 = exp_sign;
      7'b0001000: n16427 = n16329;
      7'b0000100: n16427 = exp_sign;
      7'b0000010: n16427 = n15874;
      7'b0000001: n16427 = exp_sign;
      default: n16427 = 1'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16430 = cycle_count;
      7'b0100000: n16430 = cycle_count;
      7'b0010000: n16430 = cycle_count;
      7'b0001000: n16430 = n16330;
      7'b0000100: n16430 = n16098;
      7'b0000010: n16430 = cycle_count;
      7'b0000001: n16430 = 6'b000000;
      default: n16430 = 6'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:146:17  */
  always @*
    case (n16384)
      7'b1000000: n16432 = packed_conversion_temp_mantissa;
      7'b0100000: n16432 = packed_conversion_temp_mantissa;
      7'b0010000: n16432 = packed_conversion_temp_mantissa;
      7'b0001000: n16432 = n16127;
      7'b0000100: n16432 = n16099;
      7'b0000010: n16432 = packed_conversion_temp_mantissa;
      7'b0000001: n16432 = packed_conversion_temp_mantissa;
      default: n16432 = 128'bX;
    endcase
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16507 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16508 = clkena & n16507;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16509 = n16508 ? n16432 : packed_conversion_temp_mantissa;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16510 <= n16509;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16519 = clkena ? n16411 : packed_state;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16520 <= 3'b000;
    else
      n16520 <= n16519;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16521 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16522 = clkena & n16521;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16523 = n16522 ? n16413 : bcd_digits;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16524 <= n16523;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16525 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16526 = clkena & n16525;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16527 = n16526 ? n16415 : bcd_exponent;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16528 <= n16527;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16529 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16530 = clkena & n16529;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16531 = n16530 ? n16417 : binary_mantissa;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16532 <= n16531;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16534 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16535 = clkena & n16534;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16536 = n16535 ? n16419 : decimal_exponent;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16537 <= n16536;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16538 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16539 = clkena & n16538;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16540 = n16539 ? n16421 : work_mantissa;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16541 <= n16540;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16542 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16543 = clkena & n16542;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16544 = n16543 ? n16423 : work_exponent;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16545 <= n16544;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16546 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16547 = clkena & n16546;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16548 = n16547 ? n16425 : result_sign;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16549 <= n16548;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16550 = ~n15692;
  /* TG68K_FPU_PackedDecimal.vhd:127:5  */
  assign n16551 = clkena & n16550;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16552 = n16551 ? n16427 : exp_sign;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk)
    n16553 <= n16552;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16554 = clkena ? n16430 : cycle_count;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16555 <= 6'b000000;
    else
      n16555 <= n16554;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16556 = clkena ? n16388 : n16557;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16557 <= 1'b0;
    else
      n16557 <= n16556;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16558 = clkena ? n16392 : n16559;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16559 <= 1'b0;
    else
      n16559 <= n16558;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16560 = clkena ? n16394 : n16561;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16561 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n16561 <= n16560;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16562 = clkena ? n16396 : n16563;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16563 <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n16563 <= n16562;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16564 = clkena ? n16399 : n16565;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16565 <= 1'b0;
    else
      n16565 <= n16564;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16566 = clkena ? n16403 : n16567;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16567 <= 1'b0;
    else
      n16567 <= n16566;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  assign n16568 = clkena ? n16406 : n16569;
  /* TG68K_FPU_PackedDecimal.vhd:144:9  */
  always @(posedge clk or posedge n15692)
    if (n15692)
      n16569 <= 1'b0;
    else
      n16569 <= n16568;
endmodule

module tg68k_fpu_exception_handler
  (input  clk,
   input  reset,
   input  [79:0] operation_result,
   input  operation_valid,
   input  [7:0] operation_type,
   input  [79:0] operand_a,
   input  [79:0] operand_b,
   input  overflow_flag,
   input  underflow_flag,
   input  inexact_flag,
   input  invalid_flag,
   input  divide_by_zero_flag,
   input  [31:0] fpcr,
   input  [31:0] fpsr_in,
   output [31:0] fpsr_out,
   output exception_pending,
   output [7:0] exception_vector,
   output [79:0] corrected_result);
  wire [31:0] fpsr_work;
  wire exception_detected;
  wire exception_enabled;
  wire [1:0] rounding_mode;
  wire is_nan_result;
  wire is_inf_result;
  wire is_zero_result;
  wire result_sign;
  wire [1:0] n14789;
  wire n14792;
  wire [14:0] n14793;
  wire n14795;
  wire n14796;
  wire n14797;
  wire [62:0] n14798;
  wire n14800;
  wire n14801;
  wire n14802;
  wire n14805;
  wire [14:0] n14806;
  wire n14808;
  wire n14809;
  wire n14810;
  wire [62:0] n14811;
  wire n14813;
  wire n14814;
  wire n14817;
  wire [78:0] n14818;
  wire n14820;
  wire n14823;
  wire n14860;
  wire [14:0] n14861;
  wire [30:0] n14862;
  wire [31:0] n14863;
  wire n14865;
  wire [14:0] n14866;
  wire [30:0] n14867;
  wire [31:0] n14868;
  wire n14913;
  wire n14914;
  wire n14915;
  wire [62:0] n14916;
  wire n14918;
  wire n14919;
  wire n14920;
  wire n14921;
  wire n14922;
  wire n14925;
  wire n14931;
  wire n14934;
  wire n14935;
  wire n14936;
  wire [62:0] n14937;
  wire n14939;
  wire n14940;
  wire n14941;
  wire n14942;
  wire n14943;
  wire n14946;
  wire n14952;
  wire [79:0] n14978;
  wire n14980;
  wire n14982;
  wire n14985;
  wire [15:0] n14987;
  wire [16:0] n14989;
  wire [79:0] n14991;
  wire [79:0] n14992;
  wire n14994;
  wire n14996;
  wire [15:0] n15000;
  wire [16:0] n15002;
  wire [79:0] n15004;
  wire n15006;
  wire n15008;
  wire n15009;
  wire [79:0] n15012;
  wire n15014;
  wire n15015;
  wire [79:0] n15018;
  wire n15020;
  wire [15:0] n15022;
  wire [16:0] n15024;
  wire [79:0] n15026;
  wire [2:0] n15027;
  reg [79:0] n15028;
  wire [79:0] n15029;
  wire n15031;
  wire n15033;
  wire n15036;
  wire n15037;
  wire [79:0] n15039;
  wire [79:0] n15040;
  wire n15041;
  wire n15043;
  wire n15045;
  wire n15049;
  wire n15051;
  wire n15052;
  wire n15055;
  wire [15:0] n15056;
  wire [16:0] n15057;
  wire [17:0] n15059;
  wire [61:0] n15060;
  wire [79:0] n15061;
  wire n15062;
  wire [15:0] n15063;
  wire [16:0] n15064;
  wire [17:0] n15066;
  wire [61:0] n15067;
  wire [79:0] n15068;
  wire [79:0] n15069;
  wire [79:0] n15070;
  wire n15072;
  wire n15073;
  wire n15078;
  wire n15080;
  wire n15082;
  wire n15084;
  wire [2:0] n15085;
  wire n15087;
  wire [2:0] n15089;
  localparam [7:0] n15090 = 8'b00000000;
  wire [3:0] n15092;
  wire [7:0] n15096;
  wire n15097;
  wire n15098;
  wire [7:0] n15100;
  wire n15103;
  wire n15112;
  wire n15113;
  wire n15115;
  wire n15124;
  wire [7:0] n15128;
  wire n15129;
  wire n15132;
  wire n15136;
  wire [7:0] n15138;
  wire n15139;
  wire n15143;
  wire n15144;
  wire n15145;
  wire n15148;
  wire n15149;
  wire n15150;
  wire n15153;
  wire n15154;
  wire n15155;
  wire n15159;
  wire n15160;
  wire n15161;
  wire n15165;
  wire [7:0] n15168;
  wire n15169;
  wire n15172;
  wire n15176;
  wire [7:0] n15178;
  wire n15179;
  wire n15183;
  wire n15184;
  wire n15185;
  wire n15188;
  wire n15189;
  wire n15190;
  wire n15193;
  wire n15194;
  wire n15195;
  wire n15199;
  wire n15200;
  wire n15201;
  wire n15205;
  wire [7:0] n15208;
  wire n15209;
  wire n15212;
  wire n15216;
  wire [7:0] n15218;
  wire n15219;
  wire n15223;
  wire n15224;
  wire n15225;
  wire n15228;
  wire n15229;
  wire n15230;
  wire n15233;
  wire n15234;
  wire n15235;
  wire n15239;
  wire n15240;
  wire n15241;
  wire n15245;
  wire [7:0] n15248;
  wire n15249;
  wire n15252;
  wire n15256;
  wire [7:0] n15258;
  wire n15259;
  wire n15263;
  wire n15264;
  wire n15265;
  wire n15268;
  wire n15269;
  wire n15270;
  wire n15273;
  wire n15274;
  wire n15275;
  wire n15279;
  wire n15280;
  wire n15281;
  wire n15285;
  wire [7:0] n15288;
  wire n15289;
  wire n15292;
  wire n15296;
  wire [7:0] n15298;
  wire n15299;
  wire n15303;
  wire n15304;
  wire n15305;
  wire n15308;
  wire n15309;
  wire n15310;
  wire n15313;
  wire n15314;
  wire n15315;
  wire n15319;
  wire n15320;
  wire n15321;
  wire n15325;
  wire [7:0] n15328;
  wire n15329;
  wire n15332;
  wire n15336;
  wire [7:0] n15338;
  wire n15339;
  wire n15343;
  wire n15344;
  wire n15345;
  wire n15348;
  wire n15349;
  wire n15350;
  wire n15353;
  wire n15354;
  wire n15355;
  wire n15359;
  wire n15360;
  wire n15361;
  wire n15365;
  wire [7:0] n15368;
  wire n15369;
  wire n15372;
  wire n15376;
  wire [7:0] n15378;
  wire n15379;
  wire n15384;
  wire n15385;
  wire n15389;
  wire n15390;
  wire n15394;
  wire n15395;
  wire n15400;
  wire n15401;
  wire [7:0] n15406;
  wire [7:0] n15407;
  wire [7:0] n15408;
  wire [7:0] n15411;
  wire [7:0] n15412;
  wire [7:0] n15413;
  wire [7:0] n15415;
  wire [7:0] n15416;
  wire [7:0] n15419;
  wire n15420;
  wire [7:0] n15423;
  wire n15424;
  wire n15425;
  wire [7:0] n15428;
  wire n15429;
  wire n15430;
  wire [7:0] n15433;
  wire n15434;
  wire n15435;
  wire [7:0] n15438;
  wire n15439;
  wire n15440;
  wire [7:0] n15443;
  wire n15444;
  wire n15445;
  wire [7:0] n15448;
  wire n15449;
  wire n15450;
  wire [7:0] n15453;
  wire n15454;
  wire n15455;
  wire [79:0] n15457;
  wire [31:0] n15458;
  wire [31:0] n15459;
  wire n15461;
  wire n15464;
  wire n15504;
  wire n15662;
  wire [31:0] n15663;
  reg [31:0] n15664;
  wire n15668;
  wire n15669;
  reg n15670;
  wire n15671;
  wire n15672;
  reg n15673;
  reg [31:0] n15674;
  reg n15675;
  wire [7:0] n15676;
  reg [7:0] n15677;
  reg [79:0] n15678;
  assign fpsr_out = n15674; //(module output)
  assign exception_pending = n15675; //(module output)
  assign exception_vector = n15677; //(module output)
  assign corrected_result = n15678; //(module output)
  /* TG68K_FPU_Exception_Handler.vhd:112:12  */
  assign fpsr_work = n15664; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:116:12  */
  assign exception_detected = n15670; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:117:12  */
  assign exception_enabled = n15673; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:118:12  */
  assign rounding_mode = n14789; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:122:12  */
  assign is_nan_result = n14805; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:123:12  */
  assign is_inf_result = n14817; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:124:12  */
  assign is_zero_result = n14823; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:348:17  */
  assign result_sign = n14792; // (signal)
  /* TG68K_FPU_Exception_Handler.vhd:131:26  */
  assign n14789 = fpcr[5:4]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:137:40  */
  assign n14792 = operation_result[79]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:140:28  */
  assign n14793 = operation_result[78:64]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:140:43  */
  assign n14795 = n14793 == 15'b111111111111111;
  /* TG68K_FPU_Exception_Handler.vhd:141:29  */
  assign n14796 = operation_result[63]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:141:34  */
  assign n14797 = ~n14796;
  /* TG68K_FPU_Exception_Handler.vhd:141:59  */
  assign n14798 = operation_result[62:0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:141:73  */
  assign n14800 = n14798 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Exception_Handler.vhd:141:40  */
  assign n14801 = n14797 | n14800;
  /* TG68K_FPU_Exception_Handler.vhd:140:63  */
  assign n14802 = n14801 & n14795;
  /* TG68K_FPU_Exception_Handler.vhd:140:9  */
  assign n14805 = n14802 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:148:28  */
  assign n14806 = operation_result[78:64]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:148:43  */
  assign n14808 = n14806 == 15'b111111111111111;
  /* TG68K_FPU_Exception_Handler.vhd:149:28  */
  assign n14809 = operation_result[63]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:148:63  */
  assign n14810 = n14809 & n14808;
  /* TG68K_FPU_Exception_Handler.vhd:149:59  */
  assign n14811 = operation_result[62:0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:149:73  */
  assign n14813 = n14811 == 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Exception_Handler.vhd:149:39  */
  assign n14814 = n14813 & n14810;
  /* TG68K_FPU_Exception_Handler.vhd:148:9  */
  assign n14817 = n14814 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:156:28  */
  assign n14818 = operation_result[78:0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:156:42  */
  assign n14820 = n14818 == 79'b0000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Exception_Handler.vhd:156:9  */
  assign n14823 = n14820 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:210:36  */
  assign n14860 = operand_a[79]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:211:55  */
  assign n14861 = operand_a[78:64]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:211:26  */
  assign n14862 = {16'b0, n14861};  //  uext
  /* TG68K_FPU_Exception_Handler.vhd:211:17  */
  assign n14863 = {1'b0, n14862};  //  uext
  /* TG68K_FPU_Exception_Handler.vhd:214:36  */
  assign n14865 = operand_b[79]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:215:55  */
  assign n14866 = operand_b[78:64]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:215:26  */
  assign n14867 = {16'b0, n14866};  //  uext
  /* TG68K_FPU_Exception_Handler.vhd:215:17  */
  assign n14868 = {1'b0, n14867};  //  uext
  /* TG68K_FPU_Exception_Handler.vhd:244:26  */
  assign n14913 = n14863 == 32'b00000000000000000111111111111111;
  /* TG68K_FPU_Exception_Handler.vhd:244:51  */
  assign n14914 = operand_a[63]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:244:56  */
  assign n14915 = ~n14914;
  /* TG68K_FPU_Exception_Handler.vhd:244:75  */
  assign n14916 = operand_a[62:0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:244:89  */
  assign n14918 = n14916 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Exception_Handler.vhd:244:62  */
  assign n14919 = n14915 | n14918;
  /* TG68K_FPU_Exception_Handler.vhd:244:36  */
  assign n14920 = n14919 & n14913;
  /* TG68K_FPU_Exception_Handler.vhd:246:34  */
  assign n14921 = operand_a[62]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:246:39  */
  assign n14922 = ~n14921;
  /* TG68K_FPU_Exception_Handler.vhd:246:21  */
  assign n14925 = n14922 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:244:17  */
  assign n14931 = n14920 ? n14925 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:250:26  */
  assign n14934 = n14868 == 32'b00000000000000000111111111111111;
  /* TG68K_FPU_Exception_Handler.vhd:250:51  */
  assign n14935 = operand_b[63]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:250:56  */
  assign n14936 = ~n14935;
  /* TG68K_FPU_Exception_Handler.vhd:250:75  */
  assign n14937 = operand_b[62:0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:250:89  */
  assign n14939 = n14937 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Exception_Handler.vhd:250:62  */
  assign n14940 = n14936 | n14939;
  /* TG68K_FPU_Exception_Handler.vhd:250:36  */
  assign n14941 = n14940 & n14934;
  /* TG68K_FPU_Exception_Handler.vhd:252:34  */
  assign n14942 = operand_b[62]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:252:39  */
  assign n14943 = ~n14942;
  /* TG68K_FPU_Exception_Handler.vhd:252:21  */
  assign n14946 = n14943 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:250:17  */
  assign n14952 = n14941 ? n14946 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:271:17  */
  assign n14978 = invalid_flag ? 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000 : operation_result;
  /* TG68K_FPU_Exception_Handler.vhd:271:17  */
  assign n14980 = invalid_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:271:17  */
  assign n14982 = invalid_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:282:49  */
  assign n14985 = n14860 ^ n14865;
  /* TG68K_FPU_Exception_Handler.vhd:282:61  */
  assign n14987 = {n14985, 15'b111111111111111};
  /* TG68K_FPU_Exception_Handler.vhd:282:81  */
  assign n14989 = {n14987, 1'b1};
  /* TG68K_FPU_Exception_Handler.vhd:282:87  */
  assign n14991 = {n14989, 63'b000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU_Exception_Handler.vhd:278:17  */
  assign n14992 = divide_by_zero_flag ? n14991 : n14978;
  /* TG68K_FPU_Exception_Handler.vhd:278:17  */
  assign n14994 = divide_by_zero_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:278:17  */
  assign n14996 = divide_by_zero_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:292:61  */
  assign n15000 = {result_sign, 15'b111111111111111};
  /* TG68K_FPU_Exception_Handler.vhd:292:81  */
  assign n15002 = {n15000, 1'b1};
  /* TG68K_FPU_Exception_Handler.vhd:292:87  */
  assign n15004 = {n15002, 63'b000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU_Exception_Handler.vhd:290:25  */
  assign n15006 = rounding_mode == 2'b00;
  /* TG68K_FPU_Exception_Handler.vhd:290:42  */
  assign n15008 = rounding_mode == 2'b01;
  /* TG68K_FPU_Exception_Handler.vhd:290:42  */
  assign n15009 = n15006 | n15008;
  /* TG68K_FPU_Exception_Handler.vhd:294:29  */
  assign n15012 = result_sign ? 80'b11111111111111111000000000000000000000000000000000000000000000000000000000000000 : 80'b01111111111111101111111111111111111111111111111111111111111111111111111111111111;
  /* TG68K_FPU_Exception_Handler.vhd:293:25  */
  assign n15014 = rounding_mode == 2'b10;
  /* TG68K_FPU_Exception_Handler.vhd:302:44  */
  assign n15015 = ~result_sign;
  /* TG68K_FPU_Exception_Handler.vhd:302:29  */
  assign n15018 = n15015 ? 80'b01111111111111111000000000000000000000000000000000000000000000000000000000000000 : 80'b11111111111111101111111111111111111111111111111111111111111111111111111111111111;
  /* TG68K_FPU_Exception_Handler.vhd:301:25  */
  assign n15020 = rounding_mode == 2'b11;
  /* TG68K_FPU_Exception_Handler.vhd:310:61  */
  assign n15022 = {result_sign, 15'b111111111111111};
  /* TG68K_FPU_Exception_Handler.vhd:310:81  */
  assign n15024 = {n15022, 1'b1};
  /* TG68K_FPU_Exception_Handler.vhd:310:87  */
  assign n15026 = {n15024, 63'b000000000000000000000000000000000000000000000000000000000000000};
  assign n15027 = {n15020, n15014, n15009};
  /* TG68K_FPU_Exception_Handler.vhd:289:21  */
  always @*
    case (n15027)
      3'b100: n15028 = n15018;
      3'b010: n15028 = n15012;
      3'b001: n15028 = n15004;
      default: n15028 = n15026;
    endcase
  /* TG68K_FPU_Exception_Handler.vhd:285:17  */
  assign n15029 = overflow_flag ? n15028 : n14992;
  /* TG68K_FPU_Exception_Handler.vhd:285:17  */
  assign n15031 = overflow_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:285:17  */
  assign n15033 = overflow_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:318:28  */
  assign n15036 = fpcr[11]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:318:33  */
  assign n15037 = ~n15036;
  /* TG68K_FPU_Exception_Handler.vhd:319:57  */
  assign n15039 = {result_sign, 79'b0000000000000000000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU_Exception_Handler.vhd:314:17  */
  assign n15040 = n15041 ? n15039 : n15029;
  /* TG68K_FPU_Exception_Handler.vhd:314:17  */
  assign n15041 = n15037 & underflow_flag;
  /* TG68K_FPU_Exception_Handler.vhd:314:17  */
  assign n15043 = underflow_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:314:17  */
  assign n15045 = underflow_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:324:17  */
  assign n15049 = inexact_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:324:17  */
  assign n15051 = inexact_flag ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:331:36  */
  assign n15052 = n14931 | n14952;
  /* TG68K_FPU_Exception_Handler.vhd:336:54  */
  assign n15055 = operand_a[79]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:336:70  */
  assign n15056 = operand_a[78:63]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:336:59  */
  assign n15057 = {n15055, n15056};
  /* TG68K_FPU_Exception_Handler.vhd:336:85  */
  assign n15059 = {n15057, 1'b1};
  /* TG68K_FPU_Exception_Handler.vhd:336:102  */
  assign n15060 = operand_a[61:0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:336:91  */
  assign n15061 = {n15059, n15060};
  /* TG68K_FPU_Exception_Handler.vhd:338:54  */
  assign n15062 = operand_b[79]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:338:70  */
  assign n15063 = operand_b[78:63]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:338:59  */
  assign n15064 = {n15062, n15063};
  /* TG68K_FPU_Exception_Handler.vhd:338:85  */
  assign n15066 = {n15064, 1'b1};
  /* TG68K_FPU_Exception_Handler.vhd:338:102  */
  assign n15067 = operand_b[61:0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:338:91  */
  assign n15068 = {n15066, n15067};
  /* TG68K_FPU_Exception_Handler.vhd:335:21  */
  assign n15069 = n14931 ? n15061 : n15068;
  /* TG68K_FPU_Exception_Handler.vhd:331:17  */
  assign n15070 = n15052 ? n15069 : n15040;
  /* TG68K_FPU_Exception_Handler.vhd:331:17  */
  assign n15072 = n15052 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:331:17  */
  assign n15073 = n15052 ? 1'b1 : n14982;
  /* TG68K_FPU_Exception_Handler.vhd:348:17  */
  assign n15078 = is_inf_result ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:346:17  */
  assign n15080 = is_zero_result ? 1'b0 : n15078;
  /* TG68K_FPU_Exception_Handler.vhd:346:17  */
  assign n15082 = is_zero_result ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:346:17  */
  assign n15084 = is_zero_result ? 1'b0 : result_sign;
  assign n15085 = {n15084, n15082, n15080};
  /* TG68K_FPU_Exception_Handler.vhd:344:17  */
  assign n15087 = is_nan_result ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:344:17  */
  assign n15089 = is_nan_result ? 3'b000 : n15085;
  assign n15092 = n15090[3:0]; // extract
  assign n15096 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15097 = n15096[7]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15098 = fpcr[15]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15100 = n15113 ? 8'b00110111 : n15677;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15103 = n15098 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15112 = n15098 ? 1'b0 : 1'b1;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15113 = n15098 & n15097;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15115 = n15097 ? n15103 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15124 = n15097 ? n15112 : 1'b1;
  assign n15128 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15129 = n15128[6]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15132 = fpcr[14]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15136 = n15161 ? 1'b1 : n15115;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15138 = n15160 ? 8'b00110110 : n15100;
  /* TG68K_FPU_Exception_Handler.vhd:365:29  */
  assign n15139 = n15124 & n15124;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15143 = n15165 ? 1'b0 : n15124;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15144 = n15139 & n15132;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15145 = n15124 & n15132;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15148 = n15124 & n15132;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15149 = n15144 & n15124;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15150 = n15145 & n15124;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15153 = n15148 & n15124;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15154 = n15149 & n15129;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15155 = n15150 & n15129;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15159 = n15153 & n15129;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15160 = n15154 & n15124;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15161 = n15155 & n15124;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15165 = n15159 & n15124;
  assign n15168 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15169 = n15168[5]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15172 = fpcr[13]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15176 = n15201 ? 1'b1 : n15136;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15178 = n15200 ? 8'b00110101 : n15138;
  /* TG68K_FPU_Exception_Handler.vhd:365:29  */
  assign n15179 = n15143 & n15143;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15183 = n15205 ? 1'b0 : n15143;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15184 = n15179 & n15172;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15185 = n15143 & n15172;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15188 = n15143 & n15172;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15189 = n15184 & n15143;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15190 = n15185 & n15143;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15193 = n15188 & n15143;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15194 = n15189 & n15169;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15195 = n15190 & n15169;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15199 = n15193 & n15169;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15200 = n15194 & n15143;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15201 = n15195 & n15143;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15205 = n15199 & n15143;
  assign n15208 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15209 = n15208[4]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15212 = fpcr[12]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15216 = n15241 ? 1'b1 : n15176;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15218 = n15240 ? 8'b00110100 : n15178;
  /* TG68K_FPU_Exception_Handler.vhd:365:29  */
  assign n15219 = n15183 & n15183;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15223 = n15245 ? 1'b0 : n15183;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15224 = n15219 & n15212;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15225 = n15183 & n15212;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15228 = n15183 & n15212;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15229 = n15224 & n15183;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15230 = n15225 & n15183;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15233 = n15228 & n15183;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15234 = n15229 & n15209;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15235 = n15230 & n15209;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15239 = n15233 & n15209;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15240 = n15234 & n15183;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15241 = n15235 & n15183;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15245 = n15239 & n15183;
  assign n15248 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15249 = n15248[3]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15252 = fpcr[11]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15256 = n15281 ? 1'b1 : n15216;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15258 = n15280 ? 8'b00110011 : n15218;
  /* TG68K_FPU_Exception_Handler.vhd:365:29  */
  assign n15259 = n15223 & n15223;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15263 = n15285 ? 1'b0 : n15223;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15264 = n15259 & n15252;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15265 = n15223 & n15252;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15268 = n15223 & n15252;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15269 = n15264 & n15223;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15270 = n15265 & n15223;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15273 = n15268 & n15223;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15274 = n15269 & n15249;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15275 = n15270 & n15249;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15279 = n15273 & n15249;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15280 = n15274 & n15223;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15281 = n15275 & n15223;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15285 = n15279 & n15223;
  assign n15288 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15289 = n15288[2]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15292 = fpcr[10]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15296 = n15321 ? 1'b1 : n15256;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15298 = n15320 ? 8'b00110010 : n15258;
  /* TG68K_FPU_Exception_Handler.vhd:365:29  */
  assign n15299 = n15263 & n15263;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15303 = n15325 ? 1'b0 : n15263;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15304 = n15299 & n15292;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15305 = n15263 & n15292;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15308 = n15263 & n15292;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15309 = n15304 & n15263;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15310 = n15305 & n15263;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15313 = n15308 & n15263;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15314 = n15309 & n15289;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15315 = n15310 & n15289;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15319 = n15313 & n15289;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15320 = n15314 & n15263;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15321 = n15315 & n15263;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15325 = n15319 & n15263;
  assign n15328 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15329 = n15328[1]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15332 = fpcr[9]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15336 = n15361 ? 1'b1 : n15296;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15338 = n15360 ? 8'b00110001 : n15298;
  /* TG68K_FPU_Exception_Handler.vhd:365:29  */
  assign n15339 = n15303 & n15303;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15343 = n15365 ? 1'b0 : n15303;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15344 = n15339 & n15332;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15345 = n15303 & n15332;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15348 = n15303 & n15332;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15349 = n15344 & n15303;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15350 = n15345 & n15303;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15353 = n15348 & n15303;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15354 = n15349 & n15329;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15355 = n15350 & n15329;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15359 = n15353 & n15329;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15360 = n15354 & n15303;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15361 = n15355 & n15303;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15365 = n15359 & n15303;
  assign n15368 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:358:47  */
  assign n15369 = n15368[0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:360:32  */
  assign n15372 = fpcr[8]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15376 = n15401 ? 1'b1 : n15336;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15378 = n15400 ? 8'b00110000 : n15338;
  /* TG68K_FPU_Exception_Handler.vhd:365:29  */
  assign n15379 = n15343 & n15343;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15384 = n15379 & n15372;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15385 = n15343 & n15372;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15389 = n15384 & n15343;
  /* TG68K_FPU_Exception_Handler.vhd:360:25  */
  assign n15390 = n15385 & n15343;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15394 = n15389 & n15369;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15395 = n15390 & n15369;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15400 = n15394 & n15343;
  /* TG68K_FPU_Exception_Handler.vhd:358:21  */
  assign n15401 = n15395 & n15343;
  assign n15406 = {n15089, n15087, n15092};
  /* TG68K_FPU_Exception_Handler.vhd:386:51  */
  assign n15407 = fpsr_in[23:16]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:387:50  */
  assign n15408 = fpsr_in[15:8]; // extract
  assign n15411 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:387:64  */
  assign n15412 = n15408 | n15411;
  /* TG68K_FPU_Exception_Handler.vhd:388:49  */
  assign n15413 = fpsr_in[7:0]; // extract
  assign n15415 = {n15073, n15033, n15045, n14996, n15051, 3'b000};
  /* TG68K_FPU_Exception_Handler.vhd:388:62  */
  assign n15416 = n15413 | n15415;
  assign n15419 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:390:62  */
  assign n15420 = n15419[7]; // extract
  assign n15423 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:390:92  */
  assign n15424 = n15423[6]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:390:66  */
  assign n15425 = n15420 | n15424;
  assign n15428 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:391:60  */
  assign n15429 = n15428[5]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:390:96  */
  assign n15430 = n15425 | n15429;
  assign n15433 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:391:90  */
  assign n15434 = n15433[4]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:391:64  */
  assign n15435 = n15430 | n15434;
  assign n15438 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:392:60  */
  assign n15439 = n15438[3]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:391:94  */
  assign n15440 = n15435 | n15439;
  assign n15443 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:392:90  */
  assign n15444 = n15443[2]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:392:64  */
  assign n15445 = n15440 | n15444;
  assign n15448 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:393:60  */
  assign n15449 = n15448[1]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:392:94  */
  assign n15450 = n15445 | n15449;
  assign n15453 = {1'b0, n15072, n14980, n15031, n15043, n14994, n15049, 1'b0};
  /* TG68K_FPU_Exception_Handler.vhd:393:90  */
  assign n15454 = n15453[0]; // extract
  /* TG68K_FPU_Exception_Handler.vhd:393:64  */
  assign n15455 = n15450 | n15454;
  /* TG68K_FPU_Exception_Handler.vhd:208:13  */
  assign n15457 = operation_valid ? n15070 : operation_result;
  assign n15458 = {n15406, n15407, n15412, n15416};
  /* TG68K_FPU_Exception_Handler.vhd:208:13  */
  assign n15459 = operation_valid ? n15458 : fpsr_in;
  /* TG68K_FPU_Exception_Handler.vhd:208:13  */
  assign n15461 = operation_valid ? n15455 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:208:13  */
  assign n15464 = operation_valid ? n15376 : 1'b0;
  /* TG68K_FPU_Exception_Handler.vhd:402:53  */
  assign n15504 = exception_detected & exception_enabled;
  /* TG68K_FPU_Exception_Handler.vhd:172:5  */
  assign n15662 = ~reset;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  assign n15663 = n15662 ? n15459 : fpsr_work;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  always @(posedge clk)
    n15664 <= n15663;
  /* TG68K_FPU_Exception_Handler.vhd:172:5  */
  assign n15668 = ~reset;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  assign n15669 = n15668 ? n15461 : exception_detected;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  always @(posedge clk)
    n15670 <= n15669;
  /* TG68K_FPU_Exception_Handler.vhd:172:5  */
  assign n15671 = ~reset;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  assign n15672 = n15671 ? n15464 : exception_enabled;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  always @(posedge clk)
    n15673 <= n15672;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n15674 <= 32'b00000000000000000000000000000000;
    else
      n15674 <= fpsr_work;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n15675 <= 1'b0;
    else
      n15675 <= n15504;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  assign n15676 = operation_valid ? n15378 : n15677;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n15677 <= 8'b00000000;
    else
      n15677 <= n15676;
  /* TG68K_FPU_Exception_Handler.vhd:196:9  */
  always @(posedge clk or posedge reset)
    if (reset)
      n15678 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n15678 <= n15457;
endmodule

module tg68k_fpu_movem
  (input  clk,
   input  nreset,
   input  clkena,
   input  start_movem,
   input  direction,
   input  [7:0] register_mask,
   input  predecrement,
   input  postincrement,
   input  fmovem_data_request,
   input  [2:0] fmovem_reg_index,
   input  fmovem_data_write,
   input  [79:0] fmovem_data_in,
   input  [79:0] reg_data_in,
   output movem_done,
   output movem_busy,
   output [79:0] fmovem_data_out,
   output [2:0] reg_address,
   output [79:0] reg_data_out,
   output reg_write_enable,
   output address_error);
  reg movem_state;
  wire n14671;
  wire n14675;
  wire n14678;
  wire n14684;
  wire [79:0] n14686;
  wire [2:0] n14687;
  wire [2:0] n14689;
  wire [79:0] n14690;
  wire n14693;
  wire n14694;
  wire n14696;
  wire n14698;
  wire n14700;
  wire n14704;
  wire [1:0] n14705;
  reg n14708;
  reg n14710;
  reg [79:0] n14712;
  reg [2:0] n14714;
  reg [79:0] n14716;
  reg n14719;
  reg n14722;
  reg n14724;
  wire n14761;
  reg n14762;
  wire n14765;
  reg n14766;
  wire n14767;
  reg n14768;
  wire n14769;
  wire n14770;
  wire [79:0] n14771;
  reg [79:0] n14772;
  wire n14773;
  wire n14774;
  wire [2:0] n14775;
  reg [2:0] n14776;
  wire n14777;
  wire n14778;
  wire [79:0] n14779;
  reg [79:0] n14780;
  wire n14781;
  reg n14782;
  wire n14783;
  reg n14784;
  assign movem_done = n14766; //(module output)
  assign movem_busy = n14768; //(module output)
  assign fmovem_data_out = n14772; //(module output)
  assign reg_address = n14776; //(module output)
  assign reg_data_out = n14780; //(module output)
  assign reg_write_enable = n14782; //(module output)
  assign address_error = n14784; //(module output)
  /* TG68K_FPU_MOVEM.vhd:70:16  */
  always @*
    movem_state = n14762; // (isignal)
  initial
    movem_state = 1'b0;
  /* TG68K_FPU_MOVEM.vhd:80:27  */
  assign n14671 = ~nreset;
  /* TG68K_FPU_MOVEM.vhd:98:49  */
  assign n14675 = start_movem ? 1'b1 : 1'b0;
  /* TG68K_FPU_MOVEM.vhd:98:49  */
  assign n14678 = start_movem ? 1'b1 : movem_state;
  /* TG68K_FPU_MOVEM.vhd:91:41  */
  assign n14684 = movem_state == 1'b0;
  /* TG68K_FPU_MOVEM.vhd:107:49  */
  assign n14686 = fmovem_data_request ? reg_data_in : n14772;
  /* TG68K_FPU_MOVEM.vhd:107:49  */
  assign n14687 = fmovem_data_request ? fmovem_reg_index : n14776;
  /* TG68K_FPU_MOVEM.vhd:113:49  */
  assign n14689 = fmovem_data_write ? fmovem_reg_index : n14687;
  /* TG68K_FPU_MOVEM.vhd:113:49  */
  assign n14690 = fmovem_data_write ? fmovem_data_in : n14780;
  /* TG68K_FPU_MOVEM.vhd:113:49  */
  assign n14693 = fmovem_data_write ? 1'b1 : 1'b0;
  /* TG68K_FPU_MOVEM.vhd:123:64  */
  assign n14694 = ~start_movem;
  /* TG68K_FPU_MOVEM.vhd:123:49  */
  assign n14696 = n14694 ? 1'b1 : n14766;
  /* TG68K_FPU_MOVEM.vhd:123:49  */
  assign n14698 = n14694 ? 1'b0 : n14768;
  /* TG68K_FPU_MOVEM.vhd:123:49  */
  assign n14700 = n14694 ? 1'b0 : movem_state;
  /* TG68K_FPU_MOVEM.vhd:105:41  */
  assign n14704 = movem_state == 1'b1;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14705 = {n14704, n14684};
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14708 = n14696;
      2'b01: n14708 = 1'b0;
      default: n14708 = 1'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14710 = n14698;
      2'b01: n14710 = n14675;
      default: n14710 = 1'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14712 = n14686;
      2'b01: n14712 = n14772;
      default: n14712 = 80'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14714 = n14689;
      2'b01: n14714 = n14776;
      default: n14714 = 3'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14716 = n14690;
      2'b01: n14716 = n14780;
      default: n14716 = 80'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14719 = n14693;
      2'b01: n14719 = 1'b0;
      default: n14719 = 1'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14722 = n14784;
      2'b01: n14722 = 1'b0;
      default: n14722 = 1'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:90:33  */
  always @*
    case (n14705)
      2'b10: n14724 = n14700;
      2'b01: n14724 = n14678;
      default: n14724 = 1'bX;
    endcase
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14761 = clkena ? n14724 : movem_state;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk or posedge n14671)
    if (n14671)
      n14762 <= 1'b0;
    else
      n14762 <= n14761;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14765 = clkena ? n14708 : n14766;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk or posedge n14671)
    if (n14671)
      n14766 <= 1'b0;
    else
      n14766 <= n14765;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14767 = clkena ? n14710 : n14768;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk or posedge n14671)
    if (n14671)
      n14768 <= 1'b0;
    else
      n14768 <= n14767;
  /* TG68K_FPU_MOVEM.vhd:78:9  */
  assign n14769 = ~n14671;
  /* TG68K_FPU_MOVEM.vhd:78:9  */
  assign n14770 = clkena & n14769;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14771 = n14770 ? n14712 : n14772;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk)
    n14772 <= n14771;
  /* TG68K_FPU_MOVEM.vhd:78:9  */
  assign n14773 = ~n14671;
  /* TG68K_FPU_MOVEM.vhd:78:9  */
  assign n14774 = clkena & n14773;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14775 = n14774 ? n14714 : n14776;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk)
    n14776 <= n14775;
  /* TG68K_FPU_MOVEM.vhd:78:9  */
  assign n14777 = ~n14671;
  /* TG68K_FPU_MOVEM.vhd:78:9  */
  assign n14778 = clkena & n14777;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14779 = n14778 ? n14716 : n14780;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk)
    n14780 <= n14779;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14781 = clkena ? n14719 : n14782;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk or posedge n14671)
    if (n14671)
      n14782 <= 1'b0;
    else
      n14782 <= n14781;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  assign n14783 = clkena ? n14722 : n14784;
  /* TG68K_FPU_MOVEM.vhd:88:17  */
  always @(posedge clk or posedge n14671)
    if (n14671)
      n14784 <= 1'b0;
    else
      n14784 <= n14783;
endmodule

module tg68k_fpu_constantrom
  (input  clk,
   input  nreset,
   input  [6:0] rom_offset,
   input  read_enable,
   output [79:0] constant_out,
   output constant_valid);
  wire n14575;
  wire n14578;
  wire n14580;
  wire n14582;
  wire n14584;
  wire n14586;
  wire n14588;
  wire n14590;
  wire n14592;
  wire n14594;
  wire n14596;
  wire n14598;
  wire n14600;
  wire n14602;
  wire n14604;
  wire n14606;
  wire n14608;
  wire n14610;
  wire n14612;
  wire n14614;
  wire n14616;
  wire n14618;
  wire n14620;
  wire [21:0] n14621;
  reg [79:0] n14645;
  wire n14649;
  wire [79:0] n14658;
  reg [79:0] n14659;
  reg n14660;
  assign constant_out = n14659; //(module output)
  assign constant_valid = n14660; //(module output)
  /* TG68K_FPU_ConstantROM.vhd:104:27  */
  assign n14575 = ~nreset;
  /* TG68K_FPU_ConstantROM.vhd:112:41  */
  assign n14578 = rom_offset == 7'b0000000;
  /* TG68K_FPU_ConstantROM.vhd:115:41  */
  assign n14580 = rom_offset == 7'b0001011;
  /* TG68K_FPU_ConstantROM.vhd:118:41  */
  assign n14582 = rom_offset == 7'b0001100;
  /* TG68K_FPU_ConstantROM.vhd:121:41  */
  assign n14584 = rom_offset == 7'b0001101;
  /* TG68K_FPU_ConstantROM.vhd:124:41  */
  assign n14586 = rom_offset == 7'b0001110;
  /* TG68K_FPU_ConstantROM.vhd:127:41  */
  assign n14588 = rom_offset == 7'b0001111;
  /* TG68K_FPU_ConstantROM.vhd:130:41  */
  assign n14590 = rom_offset == 7'b0110000;
  /* TG68K_FPU_ConstantROM.vhd:133:41  */
  assign n14592 = rom_offset == 7'b0110001;
  /* TG68K_FPU_ConstantROM.vhd:136:41  */
  assign n14594 = rom_offset == 7'b0110010;
  /* TG68K_FPU_ConstantROM.vhd:139:41  */
  assign n14596 = rom_offset == 7'b0110011;
  /* TG68K_FPU_ConstantROM.vhd:142:41  */
  assign n14598 = rom_offset == 7'b0110100;
  /* TG68K_FPU_ConstantROM.vhd:145:41  */
  assign n14600 = rom_offset == 7'b0110101;
  /* TG68K_FPU_ConstantROM.vhd:148:41  */
  assign n14602 = rom_offset == 7'b0110110;
  /* TG68K_FPU_ConstantROM.vhd:151:41  */
  assign n14604 = rom_offset == 7'b0110111;
  /* TG68K_FPU_ConstantROM.vhd:154:41  */
  assign n14606 = rom_offset == 7'b0111000;
  /* TG68K_FPU_ConstantROM.vhd:157:41  */
  assign n14608 = rom_offset == 7'b0111001;
  /* TG68K_FPU_ConstantROM.vhd:160:41  */
  assign n14610 = rom_offset == 7'b0111010;
  /* TG68K_FPU_ConstantROM.vhd:163:41  */
  assign n14612 = rom_offset == 7'b0111011;
  /* TG68K_FPU_ConstantROM.vhd:166:41  */
  assign n14614 = rom_offset == 7'b0111100;
  /* TG68K_FPU_ConstantROM.vhd:169:41  */
  assign n14616 = rom_offset == 7'b0111101;
  /* TG68K_FPU_ConstantROM.vhd:172:41  */
  assign n14618 = rom_offset == 7'b0111110;
  /* TG68K_FPU_ConstantROM.vhd:175:41  */
  assign n14620 = rom_offset == 7'b0111111;
  /* TG68K_FPU_Converter.vhd:303:65  */
  assign n14621 = {n14620, n14618, n14616, n14614, n14612, n14610, n14608, n14606, n14604, n14602, n14600, n14598, n14596, n14594, n14592, n14590, n14588, n14586, n14584, n14582, n14580, n14578};
  /* TG68K_FPU_ConstantROM.vhd:111:33  */
  always @*
    case (n14621)
      22'b1000000000000000000000: n14645 = 80'b01110101001001011100010001100000000100100111101010111100110010001111011010101111;
      22'b0100000000000000000000: n14645 = 80'b01011010100100101001000101111111010101000111110101110011110010000000011100000001;
      22'b0010000000000000000000: n14645 = 80'b01001101010010001100100101110110011101011000011010000001011101010000110000010111;
      22'b0001000000000000000000: n14645 = 80'b01000110101000111100011000110011010000010101110101001100000111010010001110001101;
      22'b0000100000000000000000: n14645 = 80'b01000011010100011010101001111110111010111111101110011101111110011101111010001110;
      22'b0000010000000000000000: n14645 = 80'b01000001101010001001001110111010010001111100100110000000111010011000110011100000;
      22'b0000001000000000000000: n14645 = 80'b01000000110100111000010011110000001111101001001111111111100111110100110110101010;
      22'b0000000100000000000000: n14645 = 80'b01000000011010010011101110001011010110110101000001010110111000010110101100111100;
      22'b0000000010000000000000: n14645 = 80'b01000000001101001000111000011011110010011011111100000100000000000000000000000000;
      22'b0000000001000000000000: n14645 = 80'b01000000000110011011111010111100001000000000000000000000000000000000000000000000;
      22'b0000000000100000000000: n14645 = 80'b01000000000011001001110001000000000000000000000000000000000000000000000000000000;
      22'b0000000000010000000000: n14645 = 80'b01000000000001011100100000000000000000000000000000000000000000000000000000000000;
      22'b0000000000001000000000: n14645 = 80'b01000000000000101010000000000000000000000000000000000000000000000000000000000000;
      22'b0000000000000100000000: n14645 = 80'b00111111111111111000000000000000000000000000000000000000000000000000000000000000;
      22'b0000000000000010000000: n14645 = 80'b01000000000000001001001101011101100011011101110110101010101010001010110000010111;
      22'b0000000000000001000000: n14645 = 80'b00111111111111101011000101110010000101111111011111010001110011110111100110101100;
      22'b0000000000000000100000: n14645 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
      22'b0000000000000000010000: n14645 = 80'b00111111111111011101111001011011110110001010100100110111001010000111000110010101;
      22'b0000000000000000001000: n14645 = 80'b00111111111111111011100010101010001110110010100101011100000101111111000010111100;
      22'b0000000000000000000100: n14645 = 80'b01000000000000001010110111111000010101000101100010100010101110110100101010011010;
      22'b0000000000000000000010: n14645 = 80'b00111111111111011001101000100000100110101000010011111011110011111111011110011000;
      22'b0000000000000000000001: n14645 = 80'b01000000000000001100100100001111110110101010001000100001011010001100001000110101;
      default: n14645 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU_ConstantROM.vhd:110:25  */
  assign n14649 = read_enable ? 1'b1 : 1'b0;
  /* TG68K_FPU_ConstantROM.vhd:107:17  */
  assign n14658 = read_enable ? n14645 : n14659;
  /* TG68K_FPU_ConstantROM.vhd:107:17  */
  always @(posedge clk or posedge n14575)
    if (n14575)
      n14659 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n14659 <= n14658;
  /* TG68K_FPU_ConstantROM.vhd:107:17  */
  always @(posedge clk or posedge n14575)
    if (n14575)
      n14660 <= 1'b0;
    else
      n14660 <= n14649;
endmodule

module tg68k_fpu_converter
  (input  clk,
   input  nreset,
   input  clkena,
   input  start_conversion,
   input  [2:0] source_format,
   input  [2:0] dest_format,
   input  [95:0] data_in,
   output conversion_done,
   output conversion_valid,
   output [79:0] data_out,
   output overflow,
   output underflow,
   output inexact,
   output invalid);
  reg [2:0] conv_state;
  wire dest_sign;
  wire [14:0] dest_exp;
  wire [63:0] dest_mant;
  wire [79:0] dest_extended;
  wire [31:0] int_value;
  wire [31:0] int_magnitude;
  wire [4:0] leading_zeros;
  wire single_sign;
  wire [7:0] single_exp;
  wire [22:0] single_mant;
  wire double_sign;
  wire [10:0] double_exp;
  wire [51:0] double_mant;
  wire conv_overflow;
  wire conv_underflow;
  wire conv_inexact;
  wire conv_invalid;
  wire packed_start;
  wire packed_done;
  wire packed_to_ext;
  wire [6:0] packed_k_factor;
  wire [79:0] packed_ext_out;
  wire [95:0] packed_dec_out;
  wire packed_overflow;
  wire packed_inexact;
  wire packed_invalid;
  wire \packed_converter.conversion_valid ;
  wire [15:0] n13661;
  wire [79:0] n13662;
  wire n13666;
  wire [2:0] n13669;
  wire n13671;
  wire [7:0] n13672;
  wire [31:0] n13673;
  wire n13675;
  wire [15:0] n13676;
  wire [31:0] n13677;
  wire n13679;
  wire [31:0] n13680;
  wire n13682;
  wire n13683;
  wire [7:0] n13684;
  wire [22:0] n13685;
  wire n13687;
  wire n13688;
  wire [10:0] n13689;
  wire [51:0] n13690;
  wire n13692;
  wire n13693;
  wire [14:0] n13694;
  wire [63:0] n13695;
  wire n13697;
  wire n13699;
  wire [6:0] n13700;
  reg [2:0] n13709;
  reg n13710;
  reg [14:0] n13711;
  reg [63:0] n13712;
  reg [31:0] n13713;
  reg n13714;
  reg [7:0] n13715;
  reg [22:0] n13716;
  reg n13717;
  reg [10:0] n13718;
  reg [51:0] n13719;
  reg n13721;
  reg n13723;
  reg n13725;
  reg [6:0] n13727;
  wire n13729;
  wire n13731;
  wire n13733;
  wire [31:0] n13734;
  wire n13737;
  wire [31:0] n13738;
  wire n13740;
  wire n13746;
  wire n13748;
  wire [4:0] n13751;
  wire n13755;
  wire [4:0] n13757;
  wire n13759;
  wire [4:0] n13761;
  wire n13764;
  wire n13765;
  wire [4:0] n13767;
  wire n13771;
  wire n13772;
  wire n13774;
  wire n13775;
  wire n13777;
  wire n13778;
  wire [4:0] n13780;
  wire n13784;
  wire n13785;
  wire n13787;
  wire n13788;
  wire n13790;
  wire n13791;
  wire [4:0] n13793;
  wire n13797;
  wire n13798;
  wire n13800;
  wire n13801;
  wire n13803;
  wire n13804;
  wire [4:0] n13806;
  wire n13810;
  wire n13811;
  wire n13813;
  wire n13814;
  wire n13816;
  wire n13817;
  wire [4:0] n13819;
  wire n13823;
  wire n13824;
  wire n13826;
  wire n13827;
  wire n13829;
  wire n13830;
  wire [4:0] n13832;
  wire n13836;
  wire n13837;
  wire n13839;
  wire n13840;
  wire n13842;
  wire n13843;
  wire [4:0] n13845;
  wire n13849;
  wire n13850;
  wire n13852;
  wire n13853;
  wire n13855;
  wire n13856;
  wire [4:0] n13858;
  wire n13862;
  wire n13863;
  wire n13865;
  wire n13866;
  wire n13868;
  wire n13869;
  wire [4:0] n13871;
  wire n13875;
  wire n13876;
  wire n13878;
  wire n13879;
  wire n13881;
  wire n13882;
  wire [4:0] n13884;
  wire n13888;
  wire n13889;
  wire n13891;
  wire n13892;
  wire n13894;
  wire n13895;
  wire [4:0] n13897;
  wire n13901;
  wire n13902;
  wire n13904;
  wire n13905;
  wire n13907;
  wire n13908;
  wire [4:0] n13910;
  wire n13914;
  wire n13915;
  wire n13917;
  wire n13918;
  wire n13920;
  wire n13921;
  wire [4:0] n13923;
  wire n13927;
  wire n13928;
  wire n13930;
  wire n13931;
  wire n13933;
  wire n13934;
  wire [4:0] n13936;
  wire n13940;
  wire n13941;
  wire n13943;
  wire n13944;
  wire n13946;
  wire n13947;
  wire [4:0] n13949;
  wire n13953;
  wire n13954;
  wire n13956;
  wire n13957;
  wire n13959;
  wire n13960;
  wire [4:0] n13962;
  wire n13966;
  wire n13967;
  wire n13969;
  wire n13970;
  wire n13972;
  wire n13973;
  wire [4:0] n13975;
  wire n13979;
  wire n13980;
  wire n13982;
  wire n13983;
  wire n13985;
  wire n13986;
  wire [4:0] n13988;
  wire n13992;
  wire n13993;
  wire n13995;
  wire n13996;
  wire n13998;
  wire n13999;
  wire [4:0] n14001;
  wire n14005;
  wire n14006;
  wire n14008;
  wire n14009;
  wire n14011;
  wire n14012;
  wire [4:0] n14014;
  wire n14018;
  wire n14019;
  wire n14021;
  wire n14022;
  wire n14024;
  wire n14025;
  wire [4:0] n14027;
  wire n14031;
  wire n14032;
  wire n14034;
  wire n14035;
  wire n14037;
  wire n14038;
  wire [4:0] n14040;
  wire n14044;
  wire n14045;
  wire n14047;
  wire n14048;
  wire n14050;
  wire n14051;
  wire [4:0] n14053;
  wire n14057;
  wire n14058;
  wire n14060;
  wire n14061;
  wire n14063;
  wire n14064;
  wire [4:0] n14066;
  wire n14070;
  wire n14071;
  wire n14073;
  wire n14074;
  wire n14076;
  wire n14077;
  wire [4:0] n14079;
  wire n14083;
  wire n14084;
  wire n14086;
  wire n14087;
  wire n14089;
  wire n14090;
  wire [4:0] n14092;
  wire n14096;
  wire n14097;
  wire n14099;
  wire n14100;
  wire n14102;
  wire n14103;
  wire [4:0] n14105;
  wire n14109;
  wire n14110;
  wire n14112;
  wire n14113;
  wire n14115;
  wire n14116;
  wire [4:0] n14118;
  wire n14122;
  wire n14123;
  wire n14125;
  wire n14126;
  wire n14128;
  wire n14129;
  wire [4:0] n14131;
  wire n14135;
  wire n14136;
  wire n14138;
  wire n14139;
  wire n14141;
  wire n14142;
  wire [4:0] n14144;
  wire n14149;
  wire n14152;
  wire [2:0] n14156;
  wire n14158;
  wire [14:0] n14160;
  wire [63:0] n14162;
  wire [31:0] n14163;
  wire [4:0] n14164;
  wire n14166;
  wire n14168;
  wire n14169;
  wire n14171;
  wire n14172;
  wire n14174;
  wire n14176;
  wire n14178;
  wire [23:0] n14180;
  wire [63:0] n14182;
  wire [63:0] n14184;
  wire [30:0] n14185;
  wire [31:0] n14186;
  wire [31:0] n14188;
  wire [31:0] n14190;
  wire [30:0] n14191;
  wire [14:0] n14192;
  wire [23:0] n14194;
  wire [63:0] n14196;
  wire [14:0] n14198;
  wire [63:0] n14199;
  wire [14:0] n14202;
  wire [63:0] n14204;
  wire n14207;
  wire n14209;
  wire n14211;
  wire n14213;
  wire [52:0] n14215;
  wire [63:0] n14217;
  wire [63:0] n14219;
  wire [30:0] n14220;
  wire [31:0] n14221;
  wire [31:0] n14223;
  wire [31:0] n14225;
  wire [30:0] n14226;
  wire [14:0] n14227;
  wire [52:0] n14229;
  wire [63:0] n14231;
  wire [14:0] n14233;
  wire [63:0] n14234;
  wire [14:0] n14237;
  wire [63:0] n14239;
  wire n14242;
  wire n14243;
  wire [14:0] n14244;
  wire [63:0] n14245;
  wire [2:0] n14247;
  wire n14248;
  wire [14:0] n14249;
  wire [63:0] n14250;
  wire n14251;
  wire n14252;
  wire n14253;
  wire n14255;
  wire [3:0] n14256;
  reg [2:0] n14260;
  reg n14261;
  reg [14:0] n14262;
  reg [63:0] n14263;
  reg [31:0] n14264;
  reg [4:0] n14265;
  reg n14266;
  reg n14267;
  reg n14269;
  reg n14271;
  wire n14274;
  wire n14276;
  wire [31:0] n14277;
  wire [31:0] n14279;
  wire [31:0] n14281;
  wire [30:0] n14282;
  wire [14:0] n14283;
  wire [31:0] n14284;
  wire n14286;
  wire [63:0] n14288;
  wire [31:0] n14289;
  wire n14291;
  wire [63:0] n14293;
  wire [30:0] n14294;
  wire [63:0] n14295;
  wire [63:0] n14297;
  wire [63:0] n14298;
  wire [14:0] n14300;
  wire [63:0] n14302;
  wire n14305;
  wire [15:0] n14306;
  wire [79:0] n14307;
  wire n14309;
  wire n14311;
  wire [15:0] n14312;
  wire [79:0] n14313;
  wire [1:0] n14314;
  reg n14317;
  reg n14320;
  reg [79:0] n14321;
  reg [2:0] n14325;
  reg n14327;
  reg n14329;
  reg [6:0] n14331;
  wire n14333;
  wire [79:0] n14334;
  wire n14335;
  wire n14336;
  wire n14337;
  wire n14339;
  wire n14341;
  wire [79:0] n14342;
  wire [2:0] n14344;
  wire n14345;
  wire n14346;
  wire n14347;
  wire n14349;
  wire [5:0] n14350;
  reg n14353;
  reg n14356;
  reg [79:0] n14358;
  reg [2:0] n14361;
  reg n14363;
  reg [14:0] n14365;
  reg [63:0] n14367;
  reg [31:0] n14369;
  reg [31:0] n14371;
  reg [4:0] n14373;
  reg n14375;
  reg [7:0] n14377;
  reg [22:0] n14379;
  reg n14381;
  reg [10:0] n14383;
  reg [51:0] n14385;
  reg n14388;
  reg n14391;
  reg n14394;
  reg n14397;
  reg n14400;
  reg n14402;
  reg [6:0] n14404;
  wire [2:0] n14492;
  reg [2:0] n14493;
  wire n14497;
  wire n14498;
  wire n14499;
  reg n14500;
  wire n14501;
  wire n14502;
  wire [14:0] n14503;
  reg [14:0] n14504;
  wire n14505;
  wire n14506;
  wire [63:0] n14507;
  reg [63:0] n14508;
  wire n14509;
  wire n14510;
  wire [31:0] n14511;
  reg [31:0] n14512;
  wire n14514;
  wire n14515;
  wire [31:0] n14516;
  reg [31:0] n14517;
  wire n14518;
  wire n14519;
  wire [4:0] n14520;
  reg [4:0] n14521;
  wire n14522;
  wire n14523;
  wire n14524;
  reg n14525;
  wire n14526;
  wire n14527;
  wire [7:0] n14528;
  reg [7:0] n14529;
  wire n14530;
  wire n14531;
  wire [22:0] n14532;
  reg [22:0] n14533;
  wire n14534;
  wire n14535;
  wire n14536;
  reg n14537;
  wire n14538;
  wire n14539;
  wire [10:0] n14540;
  reg [10:0] n14541;
  wire n14542;
  wire n14543;
  wire [51:0] n14544;
  reg [51:0] n14545;
  wire n14546;
  reg n14547;
  wire n14548;
  reg n14549;
  wire n14550;
  reg n14551;
  wire n14552;
  reg n14553;
  wire n14554;
  wire n14555;
  wire n14556;
  reg n14557;
  wire n14558;
  wire n14559;
  wire n14560;
  reg n14561;
  wire n14562;
  wire n14563;
  wire [6:0] n14564;
  reg [6:0] n14565;
  wire n14566;
  reg n14567;
  wire n14568;
  reg n14569;
  wire [79:0] n14570;
  reg [79:0] n14571;
  assign conversion_done = n14567; //(module output)
  assign conversion_valid = n14569; //(module output)
  assign data_out = n14571; //(module output)
  assign overflow = conv_overflow; //(module output)
  assign underflow = conv_underflow; //(module output)
  assign inexact = conv_inexact; //(module output)
  assign invalid = conv_invalid; //(module output)
  /* TG68K_FPU_Converter.vhd:82:16  */
  always @*
    conv_state = n14493; // (isignal)
  initial
    conv_state = 3'b000;
  /* TG68K_FPU_Converter.vhd:88:16  */
  assign dest_sign = n14500; // (signal)
  /* TG68K_FPU_Converter.vhd:89:16  */
  assign dest_exp = n14504; // (signal)
  /* TG68K_FPU_Converter.vhd:90:16  */
  assign dest_mant = n14508; // (signal)
  /* TG68K_FPU_Converter.vhd:91:16  */
  assign dest_extended = n13662; // (signal)
  /* TG68K_FPU_Converter.vhd:94:16  */
  assign int_value = n14512; // (signal)
  /* TG68K_FPU_Converter.vhd:96:16  */
  assign int_magnitude = n14517; // (signal)
  /* TG68K_FPU_Converter.vhd:97:16  */
  assign leading_zeros = n14521; // (signal)
  /* TG68K_FPU_Converter.vhd:100:16  */
  assign single_sign = n14525; // (signal)
  /* TG68K_FPU_Converter.vhd:101:16  */
  assign single_exp = n14529; // (signal)
  /* TG68K_FPU_Converter.vhd:102:16  */
  assign single_mant = n14533; // (signal)
  /* TG68K_FPU_Converter.vhd:105:16  */
  assign double_sign = n14537; // (signal)
  /* TG68K_FPU_Converter.vhd:106:16  */
  assign double_exp = n14541; // (signal)
  /* TG68K_FPU_Converter.vhd:107:16  */
  assign double_mant = n14545; // (signal)
  /* TG68K_FPU_Converter.vhd:110:16  */
  assign conv_overflow = n14547; // (signal)
  /* TG68K_FPU_Converter.vhd:111:16  */
  assign conv_underflow = n14549; // (signal)
  /* TG68K_FPU_Converter.vhd:112:16  */
  assign conv_inexact = n14551; // (signal)
  /* TG68K_FPU_Converter.vhd:113:16  */
  assign conv_invalid = n14553; // (signal)
  /* TG68K_FPU_Converter.vhd:116:16  */
  assign packed_start = n14557; // (signal)
  /* TG68K_FPU_Converter.vhd:119:16  */
  assign packed_to_ext = n14561; // (signal)
  /* TG68K_FPU_Converter.vhd:120:16  */
  assign packed_k_factor = n14565; // (signal)
  /* TG68K_FPU_Converter.vhd:130:9  */
  tg68k_fpu_packeddecimal packed_converter (
    .clk(clk),
    .nreset(nreset),
    .clkena(clkena),
    .start_conversion(packed_start),
    .packed_to_extended(packed_to_ext),
    .k_factor(packed_k_factor),
    .extended_in(dest_extended),
    .packed_in(data_in),
    .conversion_done(packed_done),
    .conversion_valid(),
    .extended_out(packed_ext_out),
    .packed_out(packed_dec_out),
    .overflow(packed_overflow),
    .inexact(packed_inexact),
    .invalid(packed_invalid));
  /* TG68K_FPU_Converter.vhd:158:36  */
  assign n13661 = {dest_sign, dest_exp};
  /* TG68K_FPU_Converter.vhd:158:47  */
  assign n13662 = {n13661, dest_mant};
  /* TG68K_FPU_Converter.vhd:165:27  */
  assign n13666 = ~nreset;
  /* TG68K_FPU_Converter.vhd:186:49  */
  assign n13669 = start_conversion ? 3'b001 : conv_state;
  /* TG68K_FPU_Converter.vhd:178:41  */
  assign n13671 = conv_state == 3'b000;
  /* TG68K_FPU_Converter.vhd:195:99  */
  assign n13672 = data_in[7:0]; // extract
  /* TG68K_FPU_Converter.vhd:195:78  */
  assign n13673 = {{24{n13672[7]}}, n13672}; // sext
  /* TG68K_FPU_Converter.vhd:193:57  */
  assign n13675 = source_format == 3'b110;
  /* TG68K_FPU_Converter.vhd:200:99  */
  assign n13676 = data_in[15:0]; // extract
  /* TG68K_FPU_Converter.vhd:200:78  */
  assign n13677 = {{16{n13676[15]}}, n13676}; // sext
  /* TG68K_FPU_Converter.vhd:198:57  */
  assign n13679 = source_format == 3'b100;
  /* TG68K_FPU_Converter.vhd:205:92  */
  assign n13680 = data_in[31:0]; // extract
  /* TG68K_FPU_Converter.vhd:203:57  */
  assign n13682 = source_format == 3'b000;
  /* TG68K_FPU_Converter.vhd:210:87  */
  assign n13683 = data_in[31]; // extract
  /* TG68K_FPU_Converter.vhd:211:86  */
  assign n13684 = data_in[30:23]; // extract
  /* TG68K_FPU_Converter.vhd:212:87  */
  assign n13685 = data_in[22:0]; // extract
  /* TG68K_FPU_Converter.vhd:208:57  */
  assign n13687 = source_format == 3'b001;
  /* TG68K_FPU_Converter.vhd:217:87  */
  assign n13688 = data_in[63]; // extract
  /* TG68K_FPU_Converter.vhd:218:86  */
  assign n13689 = data_in[62:52]; // extract
  /* TG68K_FPU_Converter.vhd:219:87  */
  assign n13690 = data_in[51:0]; // extract
  /* TG68K_FPU_Converter.vhd:215:57  */
  assign n13692 = source_format == 3'b101;
  /* TG68K_FPU_Converter.vhd:224:85  */
  assign n13693 = data_in[79]; // extract
  /* TG68K_FPU_Converter.vhd:225:84  */
  assign n13694 = data_in[78:64]; // extract
  /* TG68K_FPU_Converter.vhd:226:85  */
  assign n13695 = data_in[63:0]; // extract
  /* TG68K_FPU_Converter.vhd:222:57  */
  assign n13697 = source_format == 3'b010;
  /* TG68K_FPU_Converter.vhd:229:57  */
  assign n13699 = source_format == 3'b011;
  assign n13700 = {n13699, n13697, n13692, n13687, n13682, n13679, n13675};
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13709 = 3'b010;
      7'b0100000: n13709 = 3'b101;
      7'b0010000: n13709 = 3'b010;
      7'b0001000: n13709 = 3'b010;
      7'b0000100: n13709 = 3'b010;
      7'b0000010: n13709 = 3'b010;
      7'b0000001: n13709 = 3'b010;
      default: n13709 = 3'b101;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13710 = dest_sign;
      7'b0100000: n13710 = n13693;
      7'b0010000: n13710 = dest_sign;
      7'b0001000: n13710 = dest_sign;
      7'b0000100: n13710 = dest_sign;
      7'b0000010: n13710 = dest_sign;
      7'b0000001: n13710 = dest_sign;
      default: n13710 = dest_sign;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13711 = dest_exp;
      7'b0100000: n13711 = n13694;
      7'b0010000: n13711 = dest_exp;
      7'b0001000: n13711 = dest_exp;
      7'b0000100: n13711 = dest_exp;
      7'b0000010: n13711 = dest_exp;
      7'b0000001: n13711 = dest_exp;
      default: n13711 = dest_exp;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13712 = dest_mant;
      7'b0100000: n13712 = n13695;
      7'b0010000: n13712 = dest_mant;
      7'b0001000: n13712 = dest_mant;
      7'b0000100: n13712 = dest_mant;
      7'b0000010: n13712 = dest_mant;
      7'b0000001: n13712 = dest_mant;
      default: n13712 = dest_mant;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13713 = int_value;
      7'b0100000: n13713 = int_value;
      7'b0010000: n13713 = int_value;
      7'b0001000: n13713 = int_value;
      7'b0000100: n13713 = n13680;
      7'b0000010: n13713 = n13677;
      7'b0000001: n13713 = n13673;
      default: n13713 = int_value;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13714 = single_sign;
      7'b0100000: n13714 = single_sign;
      7'b0010000: n13714 = single_sign;
      7'b0001000: n13714 = n13683;
      7'b0000100: n13714 = single_sign;
      7'b0000010: n13714 = single_sign;
      7'b0000001: n13714 = single_sign;
      default: n13714 = single_sign;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13715 = single_exp;
      7'b0100000: n13715 = single_exp;
      7'b0010000: n13715 = single_exp;
      7'b0001000: n13715 = n13684;
      7'b0000100: n13715 = single_exp;
      7'b0000010: n13715 = single_exp;
      7'b0000001: n13715 = single_exp;
      default: n13715 = single_exp;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13716 = single_mant;
      7'b0100000: n13716 = single_mant;
      7'b0010000: n13716 = single_mant;
      7'b0001000: n13716 = n13685;
      7'b0000100: n13716 = single_mant;
      7'b0000010: n13716 = single_mant;
      7'b0000001: n13716 = single_mant;
      default: n13716 = single_mant;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13717 = double_sign;
      7'b0100000: n13717 = double_sign;
      7'b0010000: n13717 = n13688;
      7'b0001000: n13717 = double_sign;
      7'b0000100: n13717 = double_sign;
      7'b0000010: n13717 = double_sign;
      7'b0000001: n13717 = double_sign;
      default: n13717 = double_sign;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13718 = double_exp;
      7'b0100000: n13718 = double_exp;
      7'b0010000: n13718 = n13689;
      7'b0001000: n13718 = double_exp;
      7'b0000100: n13718 = double_exp;
      7'b0000010: n13718 = double_exp;
      7'b0000001: n13718 = double_exp;
      default: n13718 = double_exp;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13719 = double_mant;
      7'b0100000: n13719 = double_mant;
      7'b0010000: n13719 = n13690;
      7'b0001000: n13719 = double_mant;
      7'b0000100: n13719 = double_mant;
      7'b0000010: n13719 = double_mant;
      7'b0000001: n13719 = double_mant;
      default: n13719 = double_mant;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13721 = conv_invalid;
      7'b0100000: n13721 = conv_invalid;
      7'b0010000: n13721 = conv_invalid;
      7'b0001000: n13721 = conv_invalid;
      7'b0000100: n13721 = conv_invalid;
      7'b0000010: n13721 = conv_invalid;
      7'b0000001: n13721 = conv_invalid;
      default: n13721 = 1'b1;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13723 = 1'b1;
      7'b0100000: n13723 = packed_start;
      7'b0010000: n13723 = packed_start;
      7'b0001000: n13723 = packed_start;
      7'b0000100: n13723 = packed_start;
      7'b0000010: n13723 = packed_start;
      7'b0000001: n13723 = packed_start;
      default: n13723 = packed_start;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13725 = 1'b1;
      7'b0100000: n13725 = packed_to_ext;
      7'b0010000: n13725 = packed_to_ext;
      7'b0001000: n13725 = packed_to_ext;
      7'b0000100: n13725 = packed_to_ext;
      7'b0000010: n13725 = packed_to_ext;
      7'b0000001: n13725 = packed_to_ext;
      default: n13725 = packed_to_ext;
    endcase
  /* TG68K_FPU_Converter.vhd:192:49  */
  always @*
    case (n13700)
      7'b1000000: n13727 = 7'b0000000;
      7'b0100000: n13727 = packed_k_factor;
      7'b0010000: n13727 = packed_k_factor;
      7'b0001000: n13727 = packed_k_factor;
      7'b0000100: n13727 = packed_k_factor;
      7'b0000010: n13727 = packed_k_factor;
      7'b0000001: n13727 = packed_k_factor;
      default: n13727 = packed_k_factor;
    endcase
  /* TG68K_FPU_Converter.vhd:190:41  */
  assign n13729 = conv_state == 3'b001;
  /* TG68K_FPU_Converter.vhd:245:78  */
  assign n13731 = int_value == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Converter.vhd:252:86  */
  assign n13733 = $signed(int_value) < $signed(32'b00000000000000000000000000000000);
  /* TG68K_FPU_Converter.vhd:254:115  */
  assign n13734 = -int_value;
  /* TG68K_FPU_Converter.vhd:252:73  */
  assign n13737 = n13733 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Converter.vhd:252:73  */
  assign n13738 = n13733 ? n13734 : int_value;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13740 = int_magnitude[31]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13746 = n13740 ? 1'b0 : 1'b1;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13748 = int_magnitude[30]; // extract
  /* TG68K_FPU_Converter.vhd:264:89  */
  assign n13751 = n13746 ? 5'b00001 : 5'b00000;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13755 = n13764 ? 1'b0 : n13746;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13757 = n13748 ? n13751 : 5'b00000;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13759 = n13746 & n13748;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13761 = n13746 ? n13757 : 5'b00000;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13764 = n13759 & n13746;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13765 = int_magnitude[29]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13767 = n13775 ? 5'b00010 : n13761;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13771 = n13777 ? 1'b0 : n13755;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13772 = n13755 & n13765;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13774 = n13755 & n13765;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13775 = n13772 & n13755;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13777 = n13774 & n13755;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13778 = int_magnitude[28]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13780 = n13788 ? 5'b00011 : n13767;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13784 = n13790 ? 1'b0 : n13771;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13785 = n13771 & n13778;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13787 = n13771 & n13778;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13788 = n13785 & n13771;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13790 = n13787 & n13771;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13791 = int_magnitude[27]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13793 = n13801 ? 5'b00100 : n13780;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13797 = n13803 ? 1'b0 : n13784;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13798 = n13784 & n13791;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13800 = n13784 & n13791;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13801 = n13798 & n13784;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13803 = n13800 & n13784;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13804 = int_magnitude[26]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13806 = n13814 ? 5'b00101 : n13793;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13810 = n13816 ? 1'b0 : n13797;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13811 = n13797 & n13804;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13813 = n13797 & n13804;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13814 = n13811 & n13797;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13816 = n13813 & n13797;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13817 = int_magnitude[25]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13819 = n13827 ? 5'b00110 : n13806;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13823 = n13829 ? 1'b0 : n13810;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13824 = n13810 & n13817;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13826 = n13810 & n13817;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13827 = n13824 & n13810;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13829 = n13826 & n13810;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13830 = int_magnitude[24]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13832 = n13840 ? 5'b00111 : n13819;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13836 = n13842 ? 1'b0 : n13823;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13837 = n13823 & n13830;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13839 = n13823 & n13830;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13840 = n13837 & n13823;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13842 = n13839 & n13823;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13843 = int_magnitude[23]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13845 = n13853 ? 5'b01000 : n13832;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13849 = n13855 ? 1'b0 : n13836;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13850 = n13836 & n13843;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13852 = n13836 & n13843;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13853 = n13850 & n13836;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13855 = n13852 & n13836;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13856 = int_magnitude[22]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13858 = n13866 ? 5'b01001 : n13845;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13862 = n13868 ? 1'b0 : n13849;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13863 = n13849 & n13856;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13865 = n13849 & n13856;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13866 = n13863 & n13849;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13868 = n13865 & n13849;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13869 = int_magnitude[21]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13871 = n13879 ? 5'b01010 : n13858;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13875 = n13881 ? 1'b0 : n13862;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13876 = n13862 & n13869;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13878 = n13862 & n13869;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13879 = n13876 & n13862;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13881 = n13878 & n13862;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13882 = int_magnitude[20]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13884 = n13892 ? 5'b01011 : n13871;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13888 = n13894 ? 1'b0 : n13875;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13889 = n13875 & n13882;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13891 = n13875 & n13882;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13892 = n13889 & n13875;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13894 = n13891 & n13875;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13895 = int_magnitude[19]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13897 = n13905 ? 5'b01100 : n13884;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13901 = n13907 ? 1'b0 : n13888;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13902 = n13888 & n13895;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13904 = n13888 & n13895;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13905 = n13902 & n13888;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13907 = n13904 & n13888;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13908 = int_magnitude[18]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13910 = n13918 ? 5'b01101 : n13897;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13914 = n13920 ? 1'b0 : n13901;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13915 = n13901 & n13908;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13917 = n13901 & n13908;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13918 = n13915 & n13901;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13920 = n13917 & n13901;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13921 = int_magnitude[17]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13923 = n13931 ? 5'b01110 : n13910;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13927 = n13933 ? 1'b0 : n13914;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13928 = n13914 & n13921;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13930 = n13914 & n13921;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13931 = n13928 & n13914;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13933 = n13930 & n13914;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13934 = int_magnitude[16]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13936 = n13944 ? 5'b01111 : n13923;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13940 = n13946 ? 1'b0 : n13927;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13941 = n13927 & n13934;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13943 = n13927 & n13934;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13944 = n13941 & n13927;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13946 = n13943 & n13927;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13947 = int_magnitude[15]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13949 = n13957 ? 5'b10000 : n13936;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13953 = n13959 ? 1'b0 : n13940;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13954 = n13940 & n13947;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13956 = n13940 & n13947;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13957 = n13954 & n13940;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13959 = n13956 & n13940;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13960 = int_magnitude[14]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13962 = n13970 ? 5'b10001 : n13949;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13966 = n13972 ? 1'b0 : n13953;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13967 = n13953 & n13960;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13969 = n13953 & n13960;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13970 = n13967 & n13953;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13972 = n13969 & n13953;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13973 = int_magnitude[13]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13975 = n13983 ? 5'b10010 : n13962;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13979 = n13985 ? 1'b0 : n13966;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13980 = n13966 & n13973;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13982 = n13966 & n13973;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13983 = n13980 & n13966;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13985 = n13982 & n13966;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13986 = int_magnitude[12]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13988 = n13996 ? 5'b10011 : n13975;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13992 = n13998 ? 1'b0 : n13979;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13993 = n13979 & n13986;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13995 = n13979 & n13986;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13996 = n13993 & n13979;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n13998 = n13995 & n13979;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n13999 = int_magnitude[11]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14001 = n14009 ? 5'b10100 : n13988;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14005 = n14011 ? 1'b0 : n13992;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14006 = n13992 & n13999;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14008 = n13992 & n13999;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14009 = n14006 & n13992;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14011 = n14008 & n13992;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14012 = int_magnitude[10]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14014 = n14022 ? 5'b10101 : n14001;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14018 = n14024 ? 1'b0 : n14005;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14019 = n14005 & n14012;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14021 = n14005 & n14012;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14022 = n14019 & n14005;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14024 = n14021 & n14005;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14025 = int_magnitude[9]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14027 = n14035 ? 5'b10110 : n14014;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14031 = n14037 ? 1'b0 : n14018;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14032 = n14018 & n14025;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14034 = n14018 & n14025;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14035 = n14032 & n14018;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14037 = n14034 & n14018;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14038 = int_magnitude[8]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14040 = n14048 ? 5'b10111 : n14027;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14044 = n14050 ? 1'b0 : n14031;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14045 = n14031 & n14038;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14047 = n14031 & n14038;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14048 = n14045 & n14031;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14050 = n14047 & n14031;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14051 = int_magnitude[7]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14053 = n14061 ? 5'b11000 : n14040;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14057 = n14063 ? 1'b0 : n14044;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14058 = n14044 & n14051;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14060 = n14044 & n14051;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14061 = n14058 & n14044;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14063 = n14060 & n14044;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14064 = int_magnitude[6]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14066 = n14074 ? 5'b11001 : n14053;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14070 = n14076 ? 1'b0 : n14057;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14071 = n14057 & n14064;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14073 = n14057 & n14064;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14074 = n14071 & n14057;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14076 = n14073 & n14057;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14077 = int_magnitude[5]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14079 = n14087 ? 5'b11010 : n14066;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14083 = n14089 ? 1'b0 : n14070;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14084 = n14070 & n14077;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14086 = n14070 & n14077;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14087 = n14084 & n14070;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14089 = n14086 & n14070;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14090 = int_magnitude[4]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14092 = n14100 ? 5'b11011 : n14079;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14096 = n14102 ? 1'b0 : n14083;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14097 = n14083 & n14090;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14099 = n14083 & n14090;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14100 = n14097 & n14083;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14102 = n14099 & n14083;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14103 = int_magnitude[3]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14105 = n14113 ? 5'b11100 : n14092;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14109 = n14115 ? 1'b0 : n14096;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14110 = n14096 & n14103;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14112 = n14096 & n14103;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14113 = n14110 & n14096;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14115 = n14112 & n14096;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14116 = int_magnitude[2]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14118 = n14126 ? 5'b11101 : n14105;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14122 = n14128 ? 1'b0 : n14109;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14123 = n14109 & n14116;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14125 = n14109 & n14116;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14126 = n14123 & n14109;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14128 = n14125 & n14109;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14129 = int_magnitude[1]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14131 = n14139 ? 5'b11110 : n14118;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14135 = n14141 ? 1'b0 : n14122;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14136 = n14122 & n14129;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14138 = n14122 & n14129;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14139 = n14136 & n14122;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14141 = n14138 & n14122;
  /* TG68K_FPU_Converter.vhd:263:97  */
  assign n14142 = int_magnitude[0]; // extract
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14144 = n14152 ? 5'b11111 : n14131;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14149 = n14135 & n14142;
  /* TG68K_FPU_Converter.vhd:263:81  */
  assign n14152 = n14149 & n14135;
  /* TG68K_FPU_Converter.vhd:245:65  */
  assign n14156 = n13731 ? conv_state : 3'b011;
  /* TG68K_FPU_Converter.vhd:245:65  */
  assign n14158 = n13731 ? 1'b0 : n13737;
  /* TG68K_FPU_Converter.vhd:245:65  */
  assign n14160 = n13731 ? 15'b000000000000000 : dest_exp;
  /* TG68K_FPU_Converter.vhd:245:65  */
  assign n14162 = n13731 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : dest_mant;
  /* TG68K_FPU_Converter.vhd:245:65  */
  assign n14163 = n13731 ? int_magnitude : n13738;
  /* TG68K_FPU_Converter.vhd:245:65  */
  assign n14164 = n13731 ? leading_zeros : n14144;
  /* TG68K_FPU_Converter.vhd:243:57  */
  assign n14166 = source_format == 3'b110;
  /* TG68K_FPU_Converter.vhd:243:74  */
  assign n14168 = source_format == 3'b100;
  /* TG68K_FPU_Converter.vhd:243:74  */
  assign n14169 = n14166 | n14168;
  /* TG68K_FPU_Converter.vhd:243:88  */
  assign n14171 = source_format == 3'b000;
  /* TG68K_FPU_Converter.vhd:243:88  */
  assign n14172 = n14169 | n14171;
  /* TG68K_FPU_Converter.vhd:276:79  */
  assign n14174 = single_exp == 8'b00000000;
  /* TG68K_FPU_Converter.vhd:280:82  */
  assign n14176 = single_exp == 8'b11111111;
  /* TG68K_FPU_Converter.vhd:283:88  */
  assign n14178 = single_mant == 23'b00000000000000000000000;
  /* TG68K_FPU_Converter.vhd:288:98  */
  assign n14180 = {1'b1, single_mant};
  /* TG68K_FPU_Converter.vhd:288:112  */
  assign n14182 = {n14180, 40'b0000000000000000000000000000000000000000};
  /* TG68K_FPU_Converter.vhd:283:73  */
  assign n14184 = n14178 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n14182;
  /* TG68K_FPU_Converter.vhd:292:85  */
  assign n14185 = {23'b0, single_exp};  //  uext
  /* TG68K_FPU_Converter.vhd:292:118  */
  assign n14186 = {1'b0, n14185};  //  uext
  /* TG68K_FPU_Converter.vhd:292:118  */
  assign n14188 = n14186 - 32'b00000000000000000000000001111111;
  /* TG68K_FPU_Converter.vhd:292:136  */
  assign n14190 = n14188 + 32'b00000000000000000011111111111111;
  /* TG68K_FPU_Converter.vhd:293:114  */
  assign n14191 = n14190[30:0];  // trunc
  /* TG68K_FPU_Converter.vhd:293:102  */
  assign n14192 = n14191[14:0];  // trunc
  /* TG68K_FPU_Converter.vhd:295:90  */
  assign n14194 = {1'b1, single_mant};
  /* TG68K_FPU_Converter.vhd:295:104  */
  assign n14196 = {n14194, 40'b0000000000000000000000000000000000000000};
  /* TG68K_FPU_Converter.vhd:280:65  */
  assign n14198 = n14176 ? 15'b111111111111111 : n14192;
  /* TG68K_FPU_Converter.vhd:280:65  */
  assign n14199 = n14176 ? n14184 : n14196;
  /* TG68K_FPU_Converter.vhd:276:65  */
  assign n14202 = n14174 ? 15'b000000000000000 : n14198;
  /* TG68K_FPU_Converter.vhd:276:65  */
  assign n14204 = n14174 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n14199;
  /* TG68K_FPU_Converter.vhd:272:57  */
  assign n14207 = source_format == 3'b001;
  /* TG68K_FPU_Converter.vhd:303:79  */
  assign n14209 = double_exp == 11'b00000000000;
  /* TG68K_FPU_Converter.vhd:307:82  */
  assign n14211 = double_exp == 11'b11111111111;
  /* TG68K_FPU_Converter.vhd:310:88  */
  assign n14213 = double_mant == 52'b0000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Converter.vhd:315:98  */
  assign n14215 = {1'b1, double_mant};
  /* TG68K_FPU_Converter.vhd:315:112  */
  assign n14217 = {n14215, 11'b00000000000};
  /* TG68K_FPU_Converter.vhd:310:73  */
  assign n14219 = n14213 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n14217;
  /* TG68K_FPU_Converter.vhd:319:85  */
  assign n14220 = {20'b0, double_exp};  //  uext
  /* TG68K_FPU_Converter.vhd:319:118  */
  assign n14221 = {1'b0, n14220};  //  uext
  /* TG68K_FPU_Converter.vhd:319:118  */
  assign n14223 = n14221 - 32'b00000000000000000000001111111111;
  /* TG68K_FPU_Converter.vhd:319:136  */
  assign n14225 = n14223 + 32'b00000000000000000011111111111111;
  /* TG68K_FPU_Converter.vhd:320:114  */
  assign n14226 = n14225[30:0];  // trunc
  /* TG68K_FPU_Converter.vhd:320:102  */
  assign n14227 = n14226[14:0];  // trunc
  /* TG68K_FPU_Converter.vhd:322:90  */
  assign n14229 = {1'b1, double_mant};
  /* TG68K_FPU_Converter.vhd:322:104  */
  assign n14231 = {n14229, 11'b00000000000};
  /* TG68K_FPU_Converter.vhd:307:65  */
  assign n14233 = n14211 ? 15'b111111111111111 : n14227;
  /* TG68K_FPU_Converter.vhd:307:65  */
  assign n14234 = n14211 ? n14219 : n14231;
  /* TG68K_FPU_Converter.vhd:303:65  */
  assign n14237 = n14209 ? 15'b000000000000000 : n14233;
  /* TG68K_FPU_Converter.vhd:303:65  */
  assign n14239 = n14209 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n14234;
  /* TG68K_FPU_Converter.vhd:299:57  */
  assign n14242 = source_format == 3'b101;
  /* TG68K_FPU_Converter.vhd:331:100  */
  assign n14243 = packed_ext_out[79]; // extract
  /* TG68K_FPU_Converter.vhd:332:99  */
  assign n14244 = packed_ext_out[78:64]; // extract
  /* TG68K_FPU_Converter.vhd:333:100  */
  assign n14245 = packed_ext_out[63:0]; // extract
  /* TG68K_FPU_Converter.vhd:329:65  */
  assign n14247 = packed_done ? 3'b101 : conv_state;
  /* TG68K_FPU_Converter.vhd:329:65  */
  assign n14248 = packed_done ? n14243 : dest_sign;
  /* TG68K_FPU_Converter.vhd:329:65  */
  assign n14249 = packed_done ? n14244 : dest_exp;
  /* TG68K_FPU_Converter.vhd:329:65  */
  assign n14250 = packed_done ? n14245 : dest_mant;
  /* TG68K_FPU_Converter.vhd:329:65  */
  assign n14251 = packed_done ? packed_overflow : conv_overflow;
  /* TG68K_FPU_Converter.vhd:329:65  */
  assign n14252 = packed_done ? packed_inexact : conv_inexact;
  /* TG68K_FPU_Converter.vhd:329:65  */
  assign n14253 = packed_done ? packed_invalid : conv_invalid;
  /* TG68K_FPU_Converter.vhd:326:57  */
  assign n14255 = source_format == 3'b011;
  assign n14256 = {n14255, n14242, n14207, n14172};
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14260 = n14247;
      4'b0100: n14260 = 3'b101;
      4'b0010: n14260 = 3'b101;
      4'b0001: n14260 = n14156;
      default: n14260 = 3'b101;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14261 = n14248;
      4'b0100: n14261 = double_sign;
      4'b0010: n14261 = single_sign;
      4'b0001: n14261 = n14158;
      default: n14261 = dest_sign;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14262 = n14249;
      4'b0100: n14262 = n14237;
      4'b0010: n14262 = n14202;
      4'b0001: n14262 = n14160;
      default: n14262 = dest_exp;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14263 = n14250;
      4'b0100: n14263 = n14239;
      4'b0010: n14263 = n14204;
      4'b0001: n14263 = n14162;
      default: n14263 = dest_mant;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14264 = int_magnitude;
      4'b0100: n14264 = int_magnitude;
      4'b0010: n14264 = int_magnitude;
      4'b0001: n14264 = n14163;
      default: n14264 = int_magnitude;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14265 = leading_zeros;
      4'b0100: n14265 = leading_zeros;
      4'b0010: n14265 = leading_zeros;
      4'b0001: n14265 = n14164;
      default: n14265 = leading_zeros;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14266 = n14251;
      4'b0100: n14266 = conv_overflow;
      4'b0010: n14266 = conv_overflow;
      4'b0001: n14266 = conv_overflow;
      default: n14266 = conv_overflow;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14267 = n14252;
      4'b0100: n14267 = conv_inexact;
      4'b0010: n14267 = conv_inexact;
      4'b0001: n14267 = conv_inexact;
      default: n14267 = conv_inexact;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14269 = n14253;
      4'b0100: n14269 = conv_invalid;
      4'b0010: n14269 = conv_invalid;
      4'b0001: n14269 = conv_invalid;
      default: n14269 = 1'b1;
    endcase
  /* TG68K_FPU_Converter.vhd:242:49  */
  always @*
    case (n14256)
      4'b1000: n14271 = 1'b0;
      4'b0100: n14271 = packed_start;
      4'b0010: n14271 = packed_start;
      4'b0001: n14271 = packed_start;
      default: n14271 = packed_start;
    endcase
  /* TG68K_FPU_Converter.vhd:241:41  */
  assign n14274 = conv_state == 3'b010;
  /* TG68K_FPU_Converter.vhd:347:66  */
  assign n14276 = int_magnitude == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Converter.vhd:352:93  */
  assign n14277 = {27'b0, leading_zeros};  //  uext
  /* TG68K_FPU_Converter.vhd:352:93  */
  assign n14279 = 32'b00000000000000000000000000011111 - n14277;
  /* TG68K_FPU_Converter.vhd:352:87  */
  assign n14281 = 32'b00000000000000000011111111111111 + n14279;
  /* TG68K_FPU_Converter.vhd:353:98  */
  assign n14282 = n14281[30:0];  // trunc
  /* TG68K_FPU_Converter.vhd:353:86  */
  assign n14283 = n14282[14:0];  // trunc
  /* TG68K_FPU_Converter.vhd:357:74  */
  assign n14284 = {27'b0, leading_zeros};  //  uext
  /* TG68K_FPU_Converter.vhd:357:74  */
  assign n14286 = n14284 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Converter.vhd:359:92  */
  assign n14288 = {int_magnitude, 32'b00000000000000000000000000000000};
  /* TG68K_FPU_Converter.vhd:360:77  */
  assign n14289 = {27'b0, leading_zeros};  //  uext
  /* TG68K_FPU_Converter.vhd:360:77  */
  assign n14291 = $signed(n14289) <= $signed(32'b00000000000000000000000000011111);
  /* TG68K_FPU_Converter.vhd:362:129  */
  assign n14293 = {int_magnitude, 32'b00000000000000000000000000000000};
  /* TG68K_FPU_Converter.vhd:362:145  */
  assign n14294 = {26'b0, leading_zeros};  //  uext
  /* TG68K_FPU_Converter.vhd:362:95  */
  assign n14295 = n14293 << n14294;
  /* TG68K_FPU_Converter.vhd:360:57  */
  assign n14297 = n14291 ? n14295 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Converter.vhd:357:57  */
  assign n14298 = n14286 ? n14288 : n14297;
  /* TG68K_FPU_Converter.vhd:347:49  */
  assign n14300 = n14276 ? 15'b000000000000000 : n14283;
  /* TG68K_FPU_Converter.vhd:347:49  */
  assign n14302 = n14276 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n14298;
  /* TG68K_FPU_Converter.vhd:345:41  */
  assign n14305 = conv_state == 3'b011;
  /* TG68K_FPU_Converter.vhd:375:87  */
  assign n14306 = {dest_sign, dest_exp};
  /* TG68K_FPU_Converter.vhd:375:98  */
  assign n14307 = {n14306, dest_mant};
  /* TG68K_FPU_Converter.vhd:373:57  */
  assign n14309 = dest_format == 3'b010;
  /* TG68K_FPU_Converter.vhd:379:57  */
  assign n14311 = dest_format == 3'b011;
  /* TG68K_FPU_Converter.vhd:387:87  */
  assign n14312 = {dest_sign, dest_exp};
  /* TG68K_FPU_Converter.vhd:387:98  */
  assign n14313 = {n14312, dest_mant};
  assign n14314 = {n14311, n14309};
  /* TG68K_FPU_Converter.vhd:372:49  */
  always @*
    case (n14314)
      2'b10: n14317 = n14567;
      2'b01: n14317 = 1'b1;
      default: n14317 = 1'b1;
    endcase
  /* TG68K_FPU_Converter.vhd:372:49  */
  always @*
    case (n14314)
      2'b10: n14320 = n14569;
      2'b01: n14320 = 1'b1;
      default: n14320 = 1'b1;
    endcase
  /* TG68K_FPU_Converter.vhd:372:49  */
  always @*
    case (n14314)
      2'b10: n14321 = n14571;
      2'b01: n14321 = n14307;
      default: n14321 = n14313;
    endcase
  /* TG68K_FPU_Converter.vhd:372:49  */
  always @*
    case (n14314)
      2'b10: n14325 = 3'b100;
      2'b01: n14325 = 3'b000;
      default: n14325 = 3'b000;
    endcase
  /* TG68K_FPU_Converter.vhd:372:49  */
  always @*
    case (n14314)
      2'b10: n14327 = 1'b1;
      2'b01: n14327 = packed_start;
      default: n14327 = packed_start;
    endcase
  /* TG68K_FPU_Converter.vhd:372:49  */
  always @*
    case (n14314)
      2'b10: n14329 = 1'b0;
      2'b01: n14329 = packed_to_ext;
      default: n14329 = packed_to_ext;
    endcase
  /* TG68K_FPU_Converter.vhd:372:49  */
  always @*
    case (n14314)
      2'b10: n14331 = 7'b0000000;
      2'b01: n14331 = packed_k_factor;
      default: n14331 = packed_k_factor;
    endcase
  /* TG68K_FPU_Converter.vhd:370:41  */
  assign n14333 = conv_state == 3'b101;
  /* TG68K_FPU_Converter.vhd:398:83  */
  assign n14334 = packed_dec_out[79:0]; // extract
  /* TG68K_FPU_Converter.vhd:399:88  */
  assign n14335 = conv_overflow | packed_overflow;
  /* TG68K_FPU_Converter.vhd:400:86  */
  assign n14336 = conv_inexact | packed_inexact;
  /* TG68K_FPU_Converter.vhd:401:86  */
  assign n14337 = conv_invalid | packed_invalid;
  /* TG68K_FPU_Converter.vhd:396:49  */
  assign n14339 = packed_done ? 1'b1 : n14567;
  /* TG68K_FPU_Converter.vhd:396:49  */
  assign n14341 = packed_done ? 1'b1 : n14569;
  /* TG68K_FPU_Converter.vhd:396:49  */
  assign n14342 = packed_done ? n14334 : n14571;
  /* TG68K_FPU_Converter.vhd:396:49  */
  assign n14344 = packed_done ? 3'b000 : conv_state;
  /* TG68K_FPU_Converter.vhd:396:49  */
  assign n14345 = packed_done ? n14335 : conv_overflow;
  /* TG68K_FPU_Converter.vhd:396:49  */
  assign n14346 = packed_done ? n14336 : conv_inexact;
  /* TG68K_FPU_Converter.vhd:396:49  */
  assign n14347 = packed_done ? n14337 : conv_invalid;
  /* TG68K_FPU_Converter.vhd:393:41  */
  assign n14349 = conv_state == 3'b100;
  assign n14350 = {n14349, n14333, n14305, n14274, n13729, n13671};
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14353 = n14339;
      6'b010000: n14353 = n14317;
      6'b001000: n14353 = n14567;
      6'b000100: n14353 = n14567;
      6'b000010: n14353 = n14567;
      6'b000001: n14353 = 1'b0;
      default: n14353 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14356 = n14341;
      6'b010000: n14356 = n14320;
      6'b001000: n14356 = n14569;
      6'b000100: n14356 = n14569;
      6'b000010: n14356 = n14569;
      6'b000001: n14356 = 1'b0;
      default: n14356 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14358 = n14342;
      6'b010000: n14358 = n14321;
      6'b001000: n14358 = n14571;
      6'b000100: n14358 = n14571;
      6'b000010: n14358 = n14571;
      6'b000001: n14358 = n14571;
      default: n14358 = 80'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14361 = n14344;
      6'b010000: n14361 = n14325;
      6'b001000: n14361 = 3'b101;
      6'b000100: n14361 = n14260;
      6'b000010: n14361 = n13709;
      6'b000001: n14361 = n13669;
      default: n14361 = 3'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14363 = dest_sign;
      6'b010000: n14363 = dest_sign;
      6'b001000: n14363 = dest_sign;
      6'b000100: n14363 = n14261;
      6'b000010: n14363 = n13710;
      6'b000001: n14363 = dest_sign;
      default: n14363 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14365 = dest_exp;
      6'b010000: n14365 = dest_exp;
      6'b001000: n14365 = n14300;
      6'b000100: n14365 = n14262;
      6'b000010: n14365 = n13711;
      6'b000001: n14365 = dest_exp;
      default: n14365 = 15'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14367 = dest_mant;
      6'b010000: n14367 = dest_mant;
      6'b001000: n14367 = n14302;
      6'b000100: n14367 = n14263;
      6'b000010: n14367 = n13712;
      6'b000001: n14367 = dest_mant;
      default: n14367 = 64'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14369 = int_value;
      6'b010000: n14369 = int_value;
      6'b001000: n14369 = int_value;
      6'b000100: n14369 = int_value;
      6'b000010: n14369 = n13713;
      6'b000001: n14369 = int_value;
      default: n14369 = 32'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14371 = int_magnitude;
      6'b010000: n14371 = int_magnitude;
      6'b001000: n14371 = int_magnitude;
      6'b000100: n14371 = n14264;
      6'b000010: n14371 = int_magnitude;
      6'b000001: n14371 = int_magnitude;
      default: n14371 = 32'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14373 = leading_zeros;
      6'b010000: n14373 = leading_zeros;
      6'b001000: n14373 = leading_zeros;
      6'b000100: n14373 = n14265;
      6'b000010: n14373 = leading_zeros;
      6'b000001: n14373 = leading_zeros;
      default: n14373 = 5'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14375 = single_sign;
      6'b010000: n14375 = single_sign;
      6'b001000: n14375 = single_sign;
      6'b000100: n14375 = single_sign;
      6'b000010: n14375 = n13714;
      6'b000001: n14375 = single_sign;
      default: n14375 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14377 = single_exp;
      6'b010000: n14377 = single_exp;
      6'b001000: n14377 = single_exp;
      6'b000100: n14377 = single_exp;
      6'b000010: n14377 = n13715;
      6'b000001: n14377 = single_exp;
      default: n14377 = 8'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14379 = single_mant;
      6'b010000: n14379 = single_mant;
      6'b001000: n14379 = single_mant;
      6'b000100: n14379 = single_mant;
      6'b000010: n14379 = n13716;
      6'b000001: n14379 = single_mant;
      default: n14379 = 23'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14381 = double_sign;
      6'b010000: n14381 = double_sign;
      6'b001000: n14381 = double_sign;
      6'b000100: n14381 = double_sign;
      6'b000010: n14381 = n13717;
      6'b000001: n14381 = double_sign;
      default: n14381 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14383 = double_exp;
      6'b010000: n14383 = double_exp;
      6'b001000: n14383 = double_exp;
      6'b000100: n14383 = double_exp;
      6'b000010: n14383 = n13718;
      6'b000001: n14383 = double_exp;
      default: n14383 = 11'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14385 = double_mant;
      6'b010000: n14385 = double_mant;
      6'b001000: n14385 = double_mant;
      6'b000100: n14385 = double_mant;
      6'b000010: n14385 = n13719;
      6'b000001: n14385 = double_mant;
      default: n14385 = 52'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14388 = n14345;
      6'b010000: n14388 = conv_overflow;
      6'b001000: n14388 = conv_overflow;
      6'b000100: n14388 = n14266;
      6'b000010: n14388 = conv_overflow;
      6'b000001: n14388 = 1'b0;
      default: n14388 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14391 = conv_underflow;
      6'b010000: n14391 = conv_underflow;
      6'b001000: n14391 = conv_underflow;
      6'b000100: n14391 = conv_underflow;
      6'b000010: n14391 = conv_underflow;
      6'b000001: n14391 = 1'b0;
      default: n14391 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14394 = n14346;
      6'b010000: n14394 = conv_inexact;
      6'b001000: n14394 = conv_inexact;
      6'b000100: n14394 = n14267;
      6'b000010: n14394 = conv_inexact;
      6'b000001: n14394 = 1'b0;
      default: n14394 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14397 = n14347;
      6'b010000: n14397 = conv_invalid;
      6'b001000: n14397 = conv_invalid;
      6'b000100: n14397 = n14269;
      6'b000010: n14397 = n13721;
      6'b000001: n14397 = 1'b0;
      default: n14397 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14400 = 1'b0;
      6'b010000: n14400 = n14327;
      6'b001000: n14400 = packed_start;
      6'b000100: n14400 = n14271;
      6'b000010: n14400 = n13723;
      6'b000001: n14400 = packed_start;
      default: n14400 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14402 = packed_to_ext;
      6'b010000: n14402 = n14329;
      6'b001000: n14402 = packed_to_ext;
      6'b000100: n14402 = packed_to_ext;
      6'b000010: n14402 = n13725;
      6'b000001: n14402 = packed_to_ext;
      default: n14402 = 1'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:177:33  */
  always @*
    case (n14350)
      6'b100000: n14404 = packed_k_factor;
      6'b010000: n14404 = n14331;
      6'b001000: n14404 = packed_k_factor;
      6'b000100: n14404 = packed_k_factor;
      6'b000010: n14404 = n13727;
      6'b000001: n14404 = packed_k_factor;
      default: n14404 = 7'bX;
    endcase
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14492 = clkena ? n14361 : conv_state;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14493 <= 3'b000;
    else
      n14493 <= n14492;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14497 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14498 = clkena & n14497;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14499 = n14498 ? n14363 : dest_sign;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14500 <= n14499;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14501 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14502 = clkena & n14501;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14503 = n14502 ? n14365 : dest_exp;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14504 <= n14503;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14505 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14506 = clkena & n14505;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14507 = n14506 ? n14367 : dest_mant;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14508 <= n14507;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14509 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14510 = clkena & n14509;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14511 = n14510 ? n14369 : int_value;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14512 <= n14511;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14514 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14515 = clkena & n14514;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14516 = n14515 ? n14371 : int_magnitude;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14517 <= n14516;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14518 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14519 = clkena & n14518;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14520 = n14519 ? n14373 : leading_zeros;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14521 <= n14520;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14522 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14523 = clkena & n14522;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14524 = n14523 ? n14375 : single_sign;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14525 <= n14524;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14526 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14527 = clkena & n14526;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14528 = n14527 ? n14377 : single_exp;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14529 <= n14528;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14530 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14531 = clkena & n14530;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14532 = n14531 ? n14379 : single_mant;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14533 <= n14532;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14534 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14535 = clkena & n14534;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14536 = n14535 ? n14381 : double_sign;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14537 <= n14536;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14538 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14539 = clkena & n14538;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14540 = n14539 ? n14383 : double_exp;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14541 <= n14540;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14542 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14543 = clkena & n14542;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14544 = n14543 ? n14385 : double_mant;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14545 <= n14544;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14546 = clkena ? n14388 : conv_overflow;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14547 <= 1'b0;
    else
      n14547 <= n14546;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14548 = clkena ? n14391 : conv_underflow;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14549 <= 1'b0;
    else
      n14549 <= n14548;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14550 = clkena ? n14394 : conv_inexact;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14551 <= 1'b0;
    else
      n14551 <= n14550;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14552 = clkena ? n14397 : conv_invalid;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14553 <= 1'b0;
    else
      n14553 <= n14552;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14554 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14555 = clkena & n14554;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14556 = n14555 ? n14400 : packed_start;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14557 <= n14556;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14558 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14559 = clkena & n14558;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14560 = n14559 ? n14402 : packed_to_ext;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14561 <= n14560;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14562 = ~n13666;
  /* TG68K_FPU_Converter.vhd:161:9  */
  assign n14563 = clkena & n14562;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14564 = n14563 ? n14404 : packed_k_factor;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk)
    n14565 <= n14564;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14566 = clkena ? n14353 : n14567;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14567 <= 1'b0;
    else
      n14567 <= n14566;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14568 = clkena ? n14356 : n14569;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14569 <= 1'b0;
    else
      n14569 <= n14568;
  /* TG68K_FPU_Converter.vhd:175:17  */
  assign n14570 = clkena ? n14358 : n14571;
  /* TG68K_FPU_Converter.vhd:175:17  */
  always @(posedge clk or posedge n13666)
    if (n13666)
      n14571 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n14571 <= n14570;
endmodule

module tg68k_fpu_transcendental
  (input  clk,
   input  nreset,
   input  clkena,
   input  start_operation,
   input  [6:0] operation_code,
   input  [79:0] operand,
   output [79:0] result,
   output result_valid,
   output overflow,
   output underflow,
   output inexact,
   output invalid,
   output operation_busy,
   output operation_done);
  reg [2:0] trans_state;
  wire [63:0] cordic_x;
  wire [63:0] cordic_y;
  wire [63:0] cordic_z;
  wire [4:0] cordic_iteration;
  wire cordic_mode;
  wire input_sign;
  wire [14:0] input_exp;
  wire [63:0] input_mant;
  wire input_zero;
  wire input_inf;
  wire input_nan;
  wire result_sign;
  wire [14:0] result_exp;
  wire [63:0] result_mant;
  wire [79:0] series_term;
  wire [79:0] series_sum;
  wire [3:0] iteration_count;
  wire trans_overflow;
  wire trans_underflow;
  wire trans_inexact;
  wire trans_invalid;
  wire [79:0] exp_argument;
  wire [79:0] log_argument;
  wire [127:0] x_squared;
  wire [127:0] x_cubed;
  wire [127:0] x_fifth;
  wire [63:0] x3_div6;
  wire [63:0] cordic_shift_x;
  wire [63:0] cordic_shift_y;
  wire [63:0] cordic_atan_val;
  wire [63:0] x5_div120;
  wire [63:0] x_n;
  wire [63:0] a_div_x_n;
  wire [63:0] x_next;
  wire [63:0] final_mant;
  wire n11071;
  wire [14:0] n11072;
  wire [63:0] n11073;
  wire [14:0] n11074;
  wire n11076;
  wire [63:0] n11077;
  wire n11079;
  wire n11080;
  wire n11083;
  wire [14:0] n11084;
  wire n11086;
  wire n11087;
  wire n11088;
  wire [62:0] n11089;
  wire n11091;
  wire n11092;
  wire n11095;
  wire [14:0] n11096;
  wire n11098;
  wire n11099;
  wire [62:0] n11100;
  wire n11102;
  wire n11103;
  wire n11104;
  wire n11105;
  wire n11108;
  wire n11111;
  wire n11115;
  wire [2:0] n11118;
  wire [3:0] n11122;
  wire n11124;
  wire n11126;
  wire n11128;
  wire n11129;
  wire n11131;
  wire n11132;
  wire n11133;
  wire [63:0] n11136;
  wire n11138;
  wire n11140;
  wire [1:0] n11141;
  reg n11144;
  reg [14:0] n11147;
  reg [63:0] n11149;
  reg n11151;
  wire [2:0] n11154;
  wire n11155;
  wire [14:0] n11156;
  wire [63:0] n11157;
  wire n11158;
  wire [2:0] n11160;
  wire n11161;
  wire [14:0] n11163;
  wire [63:0] n11164;
  wire n11165;
  wire n11167;
  wire n11168;
  wire n11169;
  wire [2:0] n11172;
  wire n11173;
  wire [14:0] n11175;
  wire [63:0] n11177;
  wire [2:0] n11179;
  wire n11181;
  wire [14:0] n11183;
  wire [63:0] n11185;
  wire n11187;
  wire n11189;
  wire n11191;
  wire n11193;
  wire n11194;
  wire n11196;
  wire [14:0] n11199;
  wire [63:0] n11202;
  wire [2:0] n11205;
  wire n11206;
  wire [14:0] n11207;
  wire [63:0] n11208;
  wire n11211;
  wire n11213;
  wire n11214;
  wire n11216;
  wire n11217;
  wire [2:0] n11220;
  wire n11222;
  wire [14:0] n11224;
  wire [63:0] n11226;
  wire [79:0] n11227;
  wire [2:0] n11229;
  wire n11231;
  wire [14:0] n11233;
  wire [63:0] n11235;
  wire n11237;
  wire [79:0] n11238;
  wire n11240;
  wire n11242;
  wire n11243;
  wire n11245;
  wire n11246;
  wire [2:0] n11247;
  reg [2:0] n11249;
  reg n11250;
  reg [14:0] n11251;
  reg [63:0] n11252;
  reg n11253;
  reg [79:0] n11255;
  wire n11257;
  wire [31:0] n11258;
  wire n11260;
  wire n11261;
  wire n11262;
  wire [14:0] n11264;
  wire [14:0] n11266;
  wire [14:0] n11268;
  wire [14:0] n11270;
  wire [14:0] n11272;
  wire [14:0] n11274;
  wire [14:0] n11276;
  wire [14:0] n11277;
  wire [31:0] n11278;
  wire [31:0] n11280;
  wire [3:0] n11281;
  wire [31:0] n11282;
  wire n11284;
  wire [15:0] n11285;
  wire n11287;
  wire [15:0] n11288;
  wire [31:0] n11289;
  wire [31:0] n11291;
  wire [15:0] n11292;
  wire [31:0] n11293;
  wire [31:0] n11294;
  wire [63:0] n11295;
  wire [63:0] n11296;
  wire [63:0] n11297;
  wire [63:0] n11299;
  wire [31:0] n11300;
  wire [31:0] n11302;
  wire [3:0] n11303;
  wire n11304;
  wire [63:0] n11306;
  wire [63:0] n11307;
  wire [63:0] n11309;
  wire [63:0] n11310;
  wire [63:0] n11312;
  wire [63:0] n11313;
  wire [63:0] n11314;
  wire n11315;
  wire n11316;
  wire [62:0] n11317;
  wire [63:0] n11319;
  wire [14:0] n11321;
  wire [14:0] n11322;
  wire [63:0] n11323;
  wire [2:0] n11325;
  wire n11327;
  wire [14:0] n11328;
  wire [63:0] n11329;
  wire [3:0] n11330;
  wire n11332;
  wire [63:0] n11333;
  wire [63:0] n11334;
  wire [63:0] n11335;
  wire [63:0] n11336;
  wire [2:0] n11337;
  wire n11338;
  wire [14:0] n11339;
  wire [63:0] n11340;
  wire [3:0] n11341;
  wire n11342;
  wire [63:0] n11344;
  wire [63:0] n11345;
  wire [63:0] n11346;
  wire [63:0] n11347;
  wire n11349;
  wire n11351;
  wire [2:0] n11354;
  wire [4:0] n11356;
  wire n11357;
  wire [14:0] n11358;
  wire [63:0] n11359;
  wire n11361;
  wire n11363;
  wire [2:0] n11366;
  wire [4:0] n11368;
  wire n11370;
  wire [14:0] n11372;
  wire [63:0] n11374;
  wire n11376;
  wire [31:0] n11377;
  wire n11379;
  wire n11381;
  wire n11382;
  wire n11383;
  wire [62:0] n11384;
  wire n11386;
  wire n11387;
  wire [31:0] n11388;
  wire [31:0] n11390;
  wire [3:0] n11391;
  wire [2:0] n11393;
  wire n11395;
  wire [14:0] n11397;
  wire [63:0] n11399;
  wire [3:0] n11400;
  wire [79:0] n11401;
  wire [31:0] n11402;
  wire n11404;
  wire [31:0] n11405;
  wire n11407;
  wire n11409;
  wire [14:0] n11411;
  wire [30:0] n11412;
  wire [30:0] n11415;
  wire [79:0] n11416;
  wire [14:0] n11418;
  wire [30:0] n11419;
  wire [30:0] n11422;
  wire [30:0] n11423;
  wire [79:0] n11424;
  wire [79:0] n11425;
  wire [31:0] n11426;
  wire n11428;
  wire n11429;
  wire [62:0] n11430;
  wire [79:0] n11431;
  wire [79:0] n11432;
  wire [79:0] n11433;
  wire [79:0] n11434;
  wire n11435;
  wire n11436;
  wire [79:0] n11437;
  wire [79:0] n11438;
  wire [31:0] n11439;
  wire [31:0] n11441;
  wire [3:0] n11442;
  wire [14:0] n11443;
  wire n11445;
  wire [63:0] n11446;
  wire n11448;
  wire n11449;
  wire n11450;
  wire [14:0] n11451;
  wire [63:0] n11452;
  wire n11454;
  wire [14:0] n11456;
  wire [63:0] n11458;
  wire [2:0] n11460;
  wire n11461;
  wire [14:0] n11462;
  wire [63:0] n11463;
  wire [79:0] n11464;
  wire [79:0] n11465;
  wire [3:0] n11466;
  wire n11468;
  wire [2:0] n11469;
  wire n11470;
  wire [14:0] n11471;
  wire [63:0] n11472;
  wire [79:0] n11473;
  wire [79:0] n11474;
  wire [3:0] n11475;
  wire n11476;
  wire [79:0] n11477;
  wire n11479;
  wire [31:0] n11480;
  wire n11482;
  wire [31:0] n11483;
  wire [31:0] n11485;
  wire [3:0] n11486;
  wire n11488;
  wire [31:0] n11489;
  wire n11491;
  wire n11492;
  wire [14:0] n11494;
  wire [63:0] n11495;
  wire [14:0] n11498;
  wire [63:0] n11500;
  wire [2:0] n11502;
  wire n11504;
  wire [14:0] n11505;
  wire [63:0] n11506;
  wire [3:0] n11507;
  wire n11509;
  wire [31:0] n11510;
  wire n11512;
  wire [31:0] n11513;
  wire [31:0] n11515;
  wire [3:0] n11516;
  wire n11518;
  wire [31:0] n11519;
  wire n11521;
  wire n11522;
  wire [14:0] n11524;
  wire [63:0] n11525;
  wire [14:0] n11528;
  wire [63:0] n11530;
  wire [2:0] n11532;
  wire n11534;
  wire [14:0] n11535;
  wire [63:0] n11536;
  wire [3:0] n11537;
  wire n11539;
  wire [31:0] n11540;
  wire n11542;
  wire [31:0] n11543;
  wire [31:0] n11545;
  wire [3:0] n11546;
  wire [2:0] n11548;
  wire n11549;
  wire [14:0] n11551;
  wire [63:0] n11553;
  wire [79:0] n11554;
  wire [3:0] n11555;
  wire [31:0] n11556;
  wire n11558;
  wire [31:0] n11559;
  wire n11561;
  wire [31:0] n11562;
  wire [31:0] n11563;
  wire [63:0] n11564;
  wire [63:0] n11565;
  wire [63:0] n11566;
  wire [127:0] n11567;
  wire [31:0] n11568;
  wire n11570;
  wire [31:0] n11571;
  wire [31:0] n11572;
  wire [63:0] n11573;
  wire [63:0] n11574;
  wire [63:0] n11575;
  wire [127:0] n11576;
  wire [31:0] n11577;
  wire n11579;
  wire [31:0] n11580;
  wire [31:0] n11582;
  wire [63:0] n11583;
  wire [31:0] n11584;
  wire n11586;
  wire [79:0] n11587;
  wire [79:0] n11588;
  wire [31:0] n11589;
  wire n11591;
  wire [31:0] n11592;
  wire [31:0] n11593;
  wire [63:0] n11594;
  wire [63:0] n11595;
  wire [63:0] n11596;
  wire [127:0] n11597;
  wire [31:0] n11598;
  wire n11600;
  wire [63:0] n11601;
  wire [127:0] n11602;
  wire [127:0] n11604;
  wire [127:0] n11606;
  wire [63:0] n11607;
  wire [31:0] n11608;
  wire n11610;
  wire [79:0] n11611;
  wire [79:0] n11612;
  wire [79:0] n11613;
  wire [79:0] n11614;
  wire [63:0] n11615;
  wire [79:0] n11616;
  wire [127:0] n11617;
  wire [63:0] n11618;
  wire [79:0] n11619;
  wire [127:0] n11620;
  wire [63:0] n11621;
  wire [79:0] n11622;
  wire [127:0] n11623;
  wire [63:0] n11624;
  wire [63:0] n11625;
  wire [79:0] n11626;
  wire [127:0] n11627;
  wire [127:0] n11628;
  wire [63:0] n11629;
  wire [63:0] n11630;
  wire [79:0] n11631;
  wire [127:0] n11632;
  wire [127:0] n11633;
  wire [127:0] n11634;
  wire [63:0] n11635;
  wire [63:0] n11636;
  wire [31:0] n11637;
  wire [31:0] n11639;
  wire [3:0] n11640;
  wire [14:0] n11641;
  wire n11643;
  wire [14:0] n11644;
  wire [63:0] n11645;
  wire [14:0] n11647;
  wire [63:0] n11649;
  wire [2:0] n11651;
  wire n11652;
  wire [14:0] n11653;
  wire [63:0] n11654;
  wire [79:0] n11655;
  wire [3:0] n11656;
  wire n11658;
  wire n11659;
  wire [127:0] n11660;
  wire [127:0] n11661;
  wire [63:0] n11662;
  wire [63:0] n11663;
  wire [2:0] n11664;
  wire n11665;
  wire [14:0] n11666;
  wire [63:0] n11667;
  wire [79:0] n11668;
  wire [3:0] n11669;
  wire n11670;
  wire [127:0] n11671;
  wire [127:0] n11672;
  wire [127:0] n11673;
  wire [63:0] n11674;
  wire [63:0] n11675;
  wire n11677;
  wire [31:0] n11678;
  wire n11680;
  wire [31:0] n11681;
  wire [31:0] n11683;
  wire [3:0] n11684;
  wire [2:0] n11686;
  wire n11687;
  wire [14:0] n11689;
  wire [63:0] n11691;
  wire [79:0] n11692;
  wire [3:0] n11693;
  wire [31:0] n11694;
  wire n11696;
  wire [31:0] n11697;
  wire n11699;
  wire [31:0] n11700;
  wire [31:0] n11701;
  wire [63:0] n11702;
  wire [63:0] n11703;
  wire [63:0] n11704;
  wire [127:0] n11705;
  wire [31:0] n11706;
  wire n11708;
  wire [31:0] n11709;
  wire [31:0] n11710;
  wire [63:0] n11711;
  wire [63:0] n11712;
  wire [63:0] n11713;
  wire [127:0] n11714;
  wire [31:0] n11715;
  wire n11717;
  wire [31:0] n11718;
  wire [31:0] n11720;
  wire [63:0] n11721;
  wire [31:0] n11722;
  wire n11724;
  wire [79:0] n11725;
  wire [79:0] n11726;
  wire [31:0] n11727;
  wire n11729;
  wire [31:0] n11730;
  wire [31:0] n11731;
  wire [63:0] n11732;
  wire [63:0] n11733;
  wire [63:0] n11734;
  wire [127:0] n11735;
  wire [31:0] n11736;
  wire n11738;
  wire [63:0] n11739;
  wire [63:0] n11741;
  wire [31:0] n11742;
  wire n11744;
  wire [79:0] n11745;
  wire [79:0] n11746;
  wire [79:0] n11747;
  wire [79:0] n11748;
  wire [63:0] n11749;
  wire [79:0] n11750;
  wire [127:0] n11751;
  wire [63:0] n11752;
  wire [79:0] n11753;
  wire [127:0] n11754;
  wire [63:0] n11755;
  wire [79:0] n11756;
  wire [127:0] n11757;
  wire [63:0] n11758;
  wire [63:0] n11759;
  wire [79:0] n11760;
  wire [127:0] n11761;
  wire [127:0] n11762;
  wire [63:0] n11763;
  wire [63:0] n11764;
  wire [79:0] n11765;
  wire [127:0] n11766;
  wire [127:0] n11767;
  wire [127:0] n11768;
  wire [63:0] n11769;
  wire [63:0] n11770;
  wire [31:0] n11771;
  wire [31:0] n11773;
  wire [3:0] n11774;
  wire n11776;
  wire [14:0] n11778;
  wire [14:0] n11779;
  wire [63:0] n11780;
  wire [14:0] n11781;
  wire [63:0] n11782;
  wire [2:0] n11784;
  wire n11785;
  wire [14:0] n11786;
  wire [63:0] n11787;
  wire [79:0] n11788;
  wire [3:0] n11789;
  wire n11791;
  wire n11792;
  wire [127:0] n11793;
  wire [127:0] n11794;
  wire [63:0] n11795;
  wire [63:0] n11796;
  wire [2:0] n11797;
  wire n11798;
  wire [14:0] n11799;
  wire [63:0] n11800;
  wire [79:0] n11801;
  wire [3:0] n11802;
  wire n11803;
  wire [127:0] n11804;
  wire [127:0] n11805;
  wire [127:0] n11806;
  wire [63:0] n11807;
  wire [63:0] n11808;
  wire n11810;
  wire [31:0] n11811;
  wire n11813;
  wire [31:0] n11814;
  wire [31:0] n11816;
  wire [3:0] n11817;
  wire [2:0] n11819;
  wire n11821;
  wire [14:0] n11823;
  wire [63:0] n11825;
  wire [79:0] n11827;
  wire [3:0] n11828;
  wire [31:0] n11829;
  wire n11831;
  wire [31:0] n11832;
  wire n11834;
  wire [31:0] n11835;
  wire [31:0] n11836;
  wire [63:0] n11837;
  wire [63:0] n11838;
  wire [63:0] n11839;
  wire [127:0] n11840;
  wire [31:0] n11841;
  wire n11843;
  wire [63:0] n11844;
  wire [63:0] n11846;
  wire [79:0] n11847;
  wire [79:0] n11848;
  wire [31:0] n11849;
  wire n11851;
  wire [31:0] n11852;
  wire [31:0] n11853;
  wire [63:0] n11854;
  wire [63:0] n11855;
  wire [63:0] n11856;
  wire [127:0] n11857;
  wire [31:0] n11858;
  wire n11860;
  wire [63:0] n11861;
  wire [63:0] n11863;
  wire [79:0] n11864;
  wire [79:0] n11865;
  wire [31:0] n11866;
  wire n11868;
  wire [31:0] n11869;
  wire [31:0] n11870;
  wire [63:0] n11871;
  wire [63:0] n11872;
  wire [63:0] n11873;
  wire [127:0] n11874;
  wire [31:0] n11875;
  wire n11877;
  wire [63:0] n11878;
  wire [63:0] n11880;
  wire [31:0] n11881;
  wire n11883;
  wire [79:0] n11884;
  wire [79:0] n11885;
  wire [79:0] n11886;
  wire [79:0] n11887;
  wire [63:0] n11888;
  wire [79:0] n11889;
  wire [127:0] n11890;
  wire [63:0] n11891;
  wire [79:0] n11892;
  wire [127:0] n11893;
  wire [63:0] n11894;
  wire [79:0] n11895;
  wire [127:0] n11896;
  wire [127:0] n11897;
  wire [63:0] n11898;
  wire [79:0] n11899;
  wire [127:0] n11900;
  wire [127:0] n11901;
  wire [63:0] n11902;
  wire [79:0] n11903;
  wire [127:0] n11904;
  wire [127:0] n11905;
  wire [127:0] n11906;
  wire [63:0] n11907;
  wire [31:0] n11908;
  wire [31:0] n11910;
  wire [3:0] n11911;
  wire n11913;
  wire [14:0] n11915;
  wire [14:0] n11916;
  wire [63:0] n11917;
  wire [14:0] n11918;
  wire [63:0] n11919;
  wire [2:0] n11921;
  wire n11923;
  wire [14:0] n11924;
  wire [63:0] n11925;
  wire [79:0] n11926;
  wire [3:0] n11927;
  wire n11929;
  wire n11930;
  wire [127:0] n11931;
  wire [127:0] n11932;
  wire [63:0] n11933;
  wire [2:0] n11934;
  wire n11935;
  wire [14:0] n11936;
  wire [63:0] n11937;
  wire [79:0] n11938;
  wire [3:0] n11939;
  wire n11940;
  wire [127:0] n11941;
  wire [127:0] n11942;
  wire [127:0] n11943;
  wire [63:0] n11944;
  wire n11946;
  wire [31:0] n11947;
  wire n11949;
  wire n11951;
  wire [31:0] n11952;
  wire [31:0] n11954;
  wire [3:0] n11955;
  wire [2:0] n11957;
  wire n11958;
  wire [14:0] n11960;
  wire [63:0] n11962;
  wire [79:0] n11963;
  wire [3:0] n11964;
  wire [2:0] n11966;
  wire n11967;
  wire [14:0] n11969;
  wire [63:0] n11971;
  wire [79:0] n11972;
  wire [3:0] n11973;
  wire [31:0] n11974;
  wire n11976;
  wire [31:0] n11977;
  wire n11979;
  wire [31:0] n11980;
  wire [31:0] n11981;
  wire [63:0] n11982;
  wire [63:0] n11983;
  wire [63:0] n11984;
  wire [127:0] n11985;
  wire [31:0] n11986;
  wire n11988;
  wire [31:0] n11989;
  wire [31:0] n11990;
  wire [63:0] n11991;
  wire [63:0] n11992;
  wire [63:0] n11993;
  wire [127:0] n11994;
  wire [31:0] n11995;
  wire n11997;
  wire [31:0] n11998;
  wire [31:0] n12000;
  wire [63:0] n12001;
  wire [31:0] n12002;
  wire n12004;
  wire [79:0] n12005;
  wire [79:0] n12006;
  wire [31:0] n12007;
  wire n12009;
  wire [31:0] n12010;
  wire [31:0] n12011;
  wire [63:0] n12012;
  wire [63:0] n12013;
  wire [63:0] n12014;
  wire [127:0] n12015;
  wire [31:0] n12016;
  wire n12018;
  wire [63:0] n12019;
  wire [127:0] n12020;
  wire [127:0] n12022;
  wire [127:0] n12024;
  wire [63:0] n12025;
  wire [31:0] n12026;
  wire n12028;
  wire [79:0] n12029;
  wire [79:0] n12030;
  wire [79:0] n12031;
  wire [79:0] n12032;
  wire [63:0] n12033;
  wire [79:0] n12034;
  wire [127:0] n12035;
  wire [63:0] n12036;
  wire [79:0] n12037;
  wire [127:0] n12038;
  wire [63:0] n12039;
  wire [79:0] n12040;
  wire [127:0] n12041;
  wire [63:0] n12042;
  wire [63:0] n12043;
  wire [79:0] n12044;
  wire [127:0] n12045;
  wire [127:0] n12046;
  wire [63:0] n12047;
  wire [63:0] n12048;
  wire [79:0] n12049;
  wire [127:0] n12050;
  wire [127:0] n12051;
  wire [127:0] n12052;
  wire [63:0] n12053;
  wire [63:0] n12054;
  wire [31:0] n12055;
  wire [31:0] n12057;
  wire [3:0] n12058;
  wire [14:0] n12059;
  wire n12061;
  wire [14:0] n12062;
  wire [63:0] n12063;
  wire [14:0] n12065;
  wire [63:0] n12067;
  wire [2:0] n12069;
  wire n12070;
  wire [14:0] n12071;
  wire [63:0] n12072;
  wire [79:0] n12073;
  wire [3:0] n12074;
  wire n12076;
  wire n12077;
  wire [127:0] n12078;
  wire [127:0] n12079;
  wire [63:0] n12080;
  wire [63:0] n12081;
  wire [2:0] n12082;
  wire n12083;
  wire [14:0] n12084;
  wire [63:0] n12085;
  wire [79:0] n12086;
  wire [3:0] n12087;
  wire n12088;
  wire [127:0] n12089;
  wire [127:0] n12090;
  wire [127:0] n12091;
  wire [63:0] n12092;
  wire [63:0] n12093;
  wire n12095;
  wire [31:0] n12096;
  wire n12098;
  wire n12100;
  wire n12102;
  wire n12104;
  wire n12105;
  wire n12106;
  wire n12108;
  wire [1:0] n12109;
  wire n12111;
  wire n12112;
  wire [31:0] n12113;
  wire [31:0] n12115;
  wire [3:0] n12116;
  wire [2:0] n12118;
  wire n12119;
  wire [14:0] n12121;
  wire [63:0] n12123;
  wire [79:0] n12124;
  wire [3:0] n12125;
  wire [2:0] n12127;
  wire n12128;
  wire [14:0] n12130;
  wire [63:0] n12132;
  wire [79:0] n12133;
  wire [3:0] n12134;
  wire [2:0] n12136;
  wire n12138;
  wire [14:0] n12140;
  wire [63:0] n12142;
  wire [79:0] n12143;
  wire [3:0] n12144;
  wire n12146;
  wire [31:0] n12147;
  wire n12149;
  wire [31:0] n12150;
  wire n12152;
  wire [31:0] n12153;
  wire [31:0] n12154;
  wire [63:0] n12155;
  wire [63:0] n12156;
  wire [63:0] n12157;
  wire [127:0] n12158;
  wire [31:0] n12159;
  wire n12161;
  wire [31:0] n12162;
  wire [31:0] n12163;
  wire [63:0] n12164;
  wire [63:0] n12165;
  wire [63:0] n12166;
  wire [127:0] n12167;
  wire [31:0] n12168;
  wire n12170;
  wire [31:0] n12171;
  wire [31:0] n12173;
  wire [63:0] n12174;
  wire [31:0] n12175;
  wire n12177;
  wire [79:0] n12178;
  wire [79:0] n12179;
  wire [31:0] n12180;
  wire n12182;
  wire [31:0] n12183;
  wire [31:0] n12184;
  wire [63:0] n12185;
  wire [63:0] n12186;
  wire [63:0] n12187;
  wire [127:0] n12188;
  wire [31:0] n12189;
  wire n12191;
  wire [63:0] n12192;
  wire [127:0] n12193;
  wire [127:0] n12195;
  wire [127:0] n12197;
  wire [63:0] n12198;
  wire [31:0] n12199;
  wire n12201;
  wire [79:0] n12202;
  wire [79:0] n12203;
  wire [79:0] n12204;
  wire [79:0] n12205;
  wire [63:0] n12206;
  wire [79:0] n12207;
  wire [127:0] n12208;
  wire [63:0] n12209;
  wire [79:0] n12210;
  wire [127:0] n12211;
  wire [63:0] n12212;
  wire [79:0] n12213;
  wire [127:0] n12214;
  wire [63:0] n12215;
  wire [63:0] n12216;
  wire [79:0] n12217;
  wire [127:0] n12218;
  wire [127:0] n12219;
  wire [63:0] n12220;
  wire [63:0] n12221;
  wire [79:0] n12222;
  wire [127:0] n12223;
  wire [127:0] n12224;
  wire [127:0] n12225;
  wire [63:0] n12226;
  wire [63:0] n12227;
  wire [31:0] n12228;
  wire [31:0] n12230;
  wire [3:0] n12231;
  wire [14:0] n12232;
  wire [63:0] n12233;
  wire [2:0] n12235;
  wire n12236;
  wire [14:0] n12237;
  wire [63:0] n12238;
  wire [79:0] n12239;
  wire [3:0] n12240;
  wire n12242;
  wire n12243;
  wire [127:0] n12244;
  wire [127:0] n12245;
  wire [63:0] n12246;
  wire [63:0] n12247;
  wire [2:0] n12248;
  wire n12249;
  wire [14:0] n12250;
  wire [63:0] n12251;
  wire [79:0] n12252;
  wire [3:0] n12253;
  wire n12254;
  wire n12255;
  wire [127:0] n12256;
  wire [127:0] n12257;
  wire [127:0] n12258;
  wire [63:0] n12259;
  wire [63:0] n12260;
  wire n12262;
  wire [31:0] n12263;
  wire n12265;
  wire n12267;
  wire n12269;
  wire n12271;
  wire n12272;
  wire n12273;
  wire n12275;
  wire [1:0] n12276;
  wire n12278;
  wire n12279;
  wire n12280;
  wire n12281;
  wire n12283;
  wire [1:0] n12284;
  wire n12286;
  wire n12287;
  wire n12288;
  wire [31:0] n12289;
  wire [31:0] n12291;
  wire [3:0] n12292;
  wire [2:0] n12294;
  wire n12296;
  wire [14:0] n12298;
  wire [63:0] n12300;
  wire [79:0] n12302;
  wire [3:0] n12303;
  wire [2:0] n12305;
  wire n12307;
  wire [14:0] n12309;
  wire [63:0] n12311;
  wire [79:0] n12312;
  wire [3:0] n12313;
  wire [2:0] n12315;
  wire n12317;
  wire [14:0] n12319;
  wire [63:0] n12321;
  wire [79:0] n12322;
  wire [3:0] n12323;
  wire [2:0] n12325;
  wire n12327;
  wire [14:0] n12329;
  wire [63:0] n12331;
  wire [79:0] n12332;
  wire [3:0] n12333;
  wire n12335;
  wire [31:0] n12336;
  wire n12338;
  wire [31:0] n12339;
  wire n12341;
  wire [31:0] n12342;
  wire [31:0] n12343;
  wire [63:0] n12344;
  wire [63:0] n12345;
  wire [63:0] n12346;
  wire [127:0] n12347;
  wire [31:0] n12348;
  wire n12350;
  wire n12351;
  wire [79:0] n12353;
  wire [79:0] n12355;
  wire [79:0] n12356;
  wire [31:0] n12357;
  wire n12359;
  wire [31:0] n12360;
  wire [31:0] n12361;
  wire [63:0] n12362;
  wire [63:0] n12363;
  wire [63:0] n12364;
  wire [127:0] n12365;
  wire [31:0] n12366;
  wire n12368;
  wire [31:0] n12369;
  wire [31:0] n12371;
  wire [63:0] n12372;
  wire [31:0] n12373;
  wire n12375;
  wire n12376;
  wire [79:0] n12377;
  wire [79:0] n12378;
  wire [79:0] n12379;
  wire [79:0] n12380;
  wire [79:0] n12381;
  wire [31:0] n12382;
  wire n12384;
  wire [31:0] n12385;
  wire [31:0] n12386;
  wire [63:0] n12387;
  wire [63:0] n12388;
  wire [63:0] n12389;
  wire [127:0] n12390;
  wire [31:0] n12391;
  wire n12393;
  wire [63:0] n12394;
  wire [127:0] n12395;
  wire [127:0] n12397;
  wire [127:0] n12399;
  wire [63:0] n12400;
  wire [63:0] n12401;
  wire [127:0] n12402;
  wire [63:0] n12403;
  wire [79:0] n12404;
  wire [127:0] n12405;
  wire [63:0] n12406;
  wire [79:0] n12407;
  wire [127:0] n12408;
  wire [63:0] n12409;
  wire [63:0] n12410;
  wire [79:0] n12411;
  wire [127:0] n12412;
  wire [127:0] n12413;
  wire [63:0] n12414;
  wire [63:0] n12415;
  wire [79:0] n12416;
  wire [127:0] n12417;
  wire [127:0] n12418;
  wire [63:0] n12419;
  wire [63:0] n12420;
  wire [79:0] n12421;
  wire [127:0] n12422;
  wire [127:0] n12423;
  wire [127:0] n12424;
  wire [63:0] n12425;
  wire [63:0] n12426;
  wire [31:0] n12427;
  wire [31:0] n12429;
  wire [3:0] n12430;
  wire [14:0] n12431;
  wire [63:0] n12432;
  wire [2:0] n12434;
  wire n12436;
  wire [14:0] n12437;
  wire [63:0] n12438;
  wire [79:0] n12439;
  wire [3:0] n12440;
  wire n12442;
  wire n12443;
  wire [127:0] n12444;
  wire [127:0] n12445;
  wire [63:0] n12446;
  wire [63:0] n12447;
  wire [2:0] n12448;
  wire n12449;
  wire [14:0] n12450;
  wire [63:0] n12451;
  wire [79:0] n12452;
  wire [3:0] n12453;
  wire n12454;
  wire n12455;
  wire [127:0] n12456;
  wire [127:0] n12457;
  wire [127:0] n12458;
  wire [63:0] n12459;
  wire [63:0] n12460;
  wire n12462;
  wire n12464;
  wire [2:0] n12467;
  wire [4:0] n12469;
  wire n12470;
  wire [14:0] n12471;
  wire [63:0] n12472;
  wire [2:0] n12474;
  wire [4:0] n12475;
  wire n12476;
  wire [14:0] n12478;
  wire [63:0] n12480;
  wire n12482;
  wire [31:0] n12483;
  wire n12485;
  wire n12487;
  wire [31:0] n12488;
  wire [31:0] n12490;
  wire [3:0] n12491;
  wire [2:0] n12493;
  wire n12494;
  wire [14:0] n12496;
  wire [63:0] n12498;
  wire [3:0] n12499;
  wire [2:0] n12501;
  wire n12503;
  wire [14:0] n12505;
  wire [63:0] n12507;
  wire [3:0] n12508;
  wire n12510;
  wire [31:0] n12511;
  wire n12513;
  wire [31:0] n12514;
  wire [31:0] n12516;
  wire [3:0] n12517;
  wire [2:0] n12519;
  wire n12520;
  wire [14:0] n12521;
  wire [63:0] n12522;
  wire [3:0] n12523;
  wire [2:0] n12524;
  wire n12525;
  wire [14:0] n12526;
  wire [63:0] n12527;
  wire [3:0] n12528;
  wire n12530;
  wire n12531;
  wire n12533;
  wire [31:0] n12534;
  wire n12536;
  wire n12538;
  wire n12539;
  wire n12540;
  wire n12542;
  wire n12543;
  wire [31:0] n12544;
  wire [31:0] n12546;
  wire [3:0] n12547;
  wire [2:0] n12549;
  wire n12551;
  wire [14:0] n12553;
  wire [63:0] n12555;
  wire [79:0] n12557;
  wire [79:0] n12559;
  wire [3:0] n12560;
  wire n12562;
  wire [79:0] n12563;
  wire [2:0] n12565;
  wire n12567;
  wire [14:0] n12569;
  wire [63:0] n12571;
  wire [79:0] n12572;
  wire [79:0] n12573;
  wire [3:0] n12574;
  wire n12575;
  wire n12577;
  wire [79:0] n12578;
  wire [2:0] n12580;
  wire n12582;
  wire [14:0] n12584;
  wire [63:0] n12586;
  wire [79:0] n12587;
  wire [79:0] n12588;
  wire [3:0] n12589;
  wire n12590;
  wire n12591;
  wire [79:0] n12592;
  wire [31:0] n12593;
  wire n12595;
  wire [31:0] n12596;
  wire n12598;
  wire [79:0] n12599;
  wire [31:0] n12600;
  wire n12602;
  wire [15:0] n12603;
  wire [15:0] n12604;
  wire [31:0] n12605;
  wire [31:0] n12606;
  wire [31:0] n12607;
  wire [31:0] n12609;
  wire [79:0] n12610;
  wire [79:0] n12611;
  wire [31:0] n12612;
  wire n12614;
  wire [15:0] n12615;
  wire [15:0] n12616;
  wire [31:0] n12617;
  wire [31:0] n12618;
  wire [31:0] n12619;
  wire [15:0] n12620;
  wire [47:0] n12621;
  wire [47:0] n12622;
  wire [47:0] n12623;
  wire [47:0] n12625;
  wire [79:0] n12626;
  wire [79:0] n12627;
  wire [31:0] n12628;
  wire n12630;
  wire [79:0] n12632;
  wire [79:0] n12633;
  wire [79:0] n12634;
  wire [79:0] n12635;
  wire [79:0] n12636;
  wire [79:0] n12637;
  wire [79:0] n12638;
  wire [79:0] n12639;
  wire [79:0] n12640;
  wire [79:0] n12641;
  wire [31:0] n12642;
  wire [31:0] n12644;
  wire [3:0] n12645;
  wire n12646;
  wire [14:0] n12647;
  wire [63:0] n12648;
  wire [2:0] n12650;
  wire n12651;
  wire [14:0] n12652;
  wire [63:0] n12653;
  wire [79:0] n12654;
  wire [79:0] n12655;
  wire [3:0] n12656;
  wire n12658;
  wire [2:0] n12659;
  wire n12660;
  wire [14:0] n12661;
  wire [63:0] n12662;
  wire [79:0] n12663;
  wire [79:0] n12664;
  wire [3:0] n12665;
  wire n12666;
  wire n12667;
  wire n12668;
  wire [79:0] n12669;
  wire n12671;
  wire [31:0] n12672;
  wire n12674;
  wire n12676;
  wire n12677;
  wire n12678;
  wire n12680;
  wire n12681;
  wire [31:0] n12682;
  wire [31:0] n12684;
  wire [3:0] n12685;
  wire [2:0] n12687;
  wire n12689;
  wire [14:0] n12691;
  wire [63:0] n12693;
  wire [79:0] n12694;
  wire [79:0] n12695;
  wire [3:0] n12696;
  wire n12698;
  wire [79:0] n12699;
  wire [2:0] n12701;
  wire n12703;
  wire [14:0] n12705;
  wire [63:0] n12707;
  wire [79:0] n12708;
  wire [79:0] n12709;
  wire [3:0] n12710;
  wire n12711;
  wire n12713;
  wire [79:0] n12714;
  wire [2:0] n12716;
  wire n12718;
  wire [14:0] n12720;
  wire [63:0] n12722;
  wire [79:0] n12723;
  wire [79:0] n12724;
  wire [3:0] n12725;
  wire n12726;
  wire n12727;
  wire [79:0] n12728;
  wire [31:0] n12729;
  wire n12731;
  wire [31:0] n12732;
  wire n12734;
  wire [15:0] n12735;
  wire [15:0] n12736;
  wire [31:0] n12737;
  wire [31:0] n12738;
  wire [31:0] n12739;
  wire [31:0] n12741;
  wire [79:0] n12742;
  wire [79:0] n12743;
  wire [31:0] n12744;
  wire n12746;
  wire [15:0] n12747;
  wire [15:0] n12748;
  wire [31:0] n12749;
  wire [31:0] n12750;
  wire [31:0] n12751;
  wire [15:0] n12752;
  wire [47:0] n12753;
  wire [47:0] n12754;
  wire [47:0] n12755;
  wire [47:0] n12757;
  wire [79:0] n12758;
  wire [79:0] n12759;
  wire [31:0] n12760;
  wire n12762;
  wire [79:0] n12764;
  wire [79:0] n12765;
  wire [79:0] n12766;
  wire [79:0] n12767;
  wire [79:0] n12768;
  wire [79:0] n12769;
  wire [79:0] n12770;
  wire [79:0] n12771;
  wire [31:0] n12772;
  wire [31:0] n12774;
  wire [3:0] n12775;
  wire n12776;
  wire [14:0] n12777;
  wire [63:0] n12778;
  wire [2:0] n12780;
  wire n12781;
  wire [14:0] n12782;
  wire [63:0] n12783;
  wire [79:0] n12784;
  wire [79:0] n12785;
  wire [3:0] n12786;
  wire n12788;
  wire [2:0] n12789;
  wire n12790;
  wire [14:0] n12791;
  wire [63:0] n12792;
  wire [79:0] n12793;
  wire [79:0] n12794;
  wire [3:0] n12795;
  wire n12796;
  wire n12797;
  wire n12798;
  wire [79:0] n12799;
  wire n12801;
  wire [31:0] n12802;
  wire n12804;
  wire n12806;
  wire n12807;
  wire n12809;
  wire n12811;
  wire n12812;
  wire n12813;
  wire [31:0] n12814;
  wire [31:0] n12816;
  wire [3:0] n12817;
  wire [2:0] n12819;
  wire n12821;
  wire [14:0] n12823;
  wire [63:0] n12825;
  wire [79:0] n12826;
  wire [79:0] n12827;
  wire [3:0] n12828;
  wire [79:0] n12829;
  wire [2:0] n12831;
  wire n12833;
  wire [14:0] n12835;
  wire [63:0] n12837;
  wire [79:0] n12838;
  wire [79:0] n12839;
  wire [3:0] n12840;
  wire [79:0] n12841;
  wire [2:0] n12843;
  wire n12845;
  wire [14:0] n12847;
  wire [63:0] n12849;
  wire [79:0] n12850;
  wire [79:0] n12851;
  wire [3:0] n12852;
  wire n12854;
  wire [79:0] n12855;
  wire [31:0] n12856;
  wire n12858;
  wire [31:0] n12859;
  wire n12861;
  wire [15:0] n12862;
  wire [15:0] n12863;
  wire [31:0] n12864;
  wire [31:0] n12865;
  wire [31:0] n12866;
  wire [31:0] n12868;
  wire [79:0] n12869;
  wire [78:0] n12871;
  wire [79:0] n12872;
  wire [31:0] n12873;
  wire n12875;
  wire [15:0] n12876;
  wire [15:0] n12877;
  wire [31:0] n12878;
  wire [31:0] n12879;
  wire [31:0] n12880;
  wire [15:0] n12881;
  wire [47:0] n12882;
  wire [47:0] n12883;
  wire [47:0] n12884;
  wire [47:0] n12886;
  wire [79:0] n12887;
  wire [79:0] n12888;
  wire [31:0] n12889;
  wire n12891;
  wire [79:0] n12893;
  wire [78:0] n12895;
  wire [79:0] n12896;
  wire [79:0] n12897;
  wire [79:0] n12898;
  wire [79:0] n12899;
  wire [79:0] n12900;
  wire [79:0] n12901;
  wire [79:0] n12902;
  wire [79:0] n12903;
  wire [79:0] n12904;
  wire [31:0] n12905;
  wire [31:0] n12907;
  wire [3:0] n12908;
  wire n12909;
  wire [14:0] n12910;
  wire [63:0] n12911;
  wire [2:0] n12913;
  wire n12914;
  wire [14:0] n12915;
  wire [63:0] n12916;
  wire [79:0] n12917;
  wire [79:0] n12918;
  wire [3:0] n12919;
  wire n12921;
  wire [2:0] n12922;
  wire n12923;
  wire [14:0] n12924;
  wire [63:0] n12925;
  wire [79:0] n12926;
  wire [79:0] n12927;
  wire [3:0] n12928;
  wire n12929;
  wire n12930;
  wire [79:0] n12931;
  wire n12933;
  wire [31:0] n12934;
  wire n12936;
  wire [31:0] n12937;
  wire [31:0] n12939;
  wire [3:0] n12940;
  wire [2:0] n12942;
  wire n12944;
  wire [14:0] n12946;
  wire [63:0] n12948;
  wire [3:0] n12949;
  wire [31:0] n12950;
  wire n12952;
  wire [31:0] n12953;
  wire [31:0] n12955;
  wire [3:0] n12956;
  wire n12958;
  wire n12959;
  wire n12960;
  wire n12962;
  wire n12963;
  wire [13:0] n12964;
  wire [14:0] n12965;
  wire [14:0] n12967;
  wire [14:0] n12969;
  wire n12971;
  wire [14:0] n12973;
  wire n12974;
  wire n12976;
  wire [2:0] n12978;
  wire n12980;
  wire [14:0] n12981;
  wire [63:0] n12983;
  wire [3:0] n12984;
  wire n12985;
  wire n12986;
  wire [2:0] n12987;
  wire n12988;
  wire [14:0] n12989;
  wire [63:0] n12990;
  wire [3:0] n12991;
  wire n12992;
  wire n12993;
  wire n12995;
  wire n12997;
  wire [31:0] n12998;
  wire n13000;
  wire [31:0] n13001;
  wire [31:0] n13003;
  wire [3:0] n13004;
  wire [2:0] n13006;
  wire n13008;
  wire [14:0] n13010;
  wire [63:0] n13012;
  wire [3:0] n13013;
  wire [31:0] n13014;
  wire n13016;
  wire [31:0] n13017;
  wire [31:0] n13019;
  wire [3:0] n13020;
  wire n13022;
  wire n13023;
  wire n13024;
  wire n13026;
  wire n13027;
  wire [14:0] n13028;
  wire [14:0] n13030;
  wire [14:0] n13032;
  wire [14:0] n13034;
  wire n13036;
  wire [14:0] n13038;
  wire n13039;
  wire n13041;
  wire [2:0] n13043;
  wire n13045;
  wire [14:0] n13046;
  wire [63:0] n13048;
  wire [3:0] n13049;
  wire n13050;
  wire n13051;
  wire [2:0] n13052;
  wire n13053;
  wire [14:0] n13054;
  wire [63:0] n13055;
  wire [3:0] n13056;
  wire n13057;
  wire n13058;
  wire n13060;
  wire n13062;
  wire [18:0] n13063;
  reg [2:0] n13065;
  reg [4:0] n13066;
  reg n13068;
  reg [14:0] n13070;
  reg [63:0] n13072;
  reg [79:0] n13073;
  reg [79:0] n13074;
  reg [3:0] n13075;
  reg n13076;
  reg n13077;
  reg n13080;
  reg n13082;
  reg [79:0] n13083;
  reg [79:0] n13084;
  reg [127:0] n13085;
  reg [127:0] n13086;
  reg [127:0] n13087;
  reg [63:0] n13088;
  reg [63:0] n13089;
  reg [63:0] n13090;
  reg [63:0] n13091;
  reg [63:0] n13092;
  reg [63:0] n13093;
  wire n13095;
  wire n13097;
  wire [31:0] n13098;
  wire n13100;
  wire [29:0] n13101;
  wire [63:0] n13102;
  wire [31:0] n13103;
  wire [31:0] n13105;
  wire [4:0] n13106;
  wire n13108;
  wire n13110;
  wire n13111;
  wire [29:0] n13112;
  wire [63:0] n13113;
  wire [29:0] n13114;
  wire [63:0] n13115;
  wire [31:0] n13116;
  wire [31:0] n13118;
  wire [4:0] n13119;
  wire n13121;
  wire [1:0] n13122;
  reg [2:0] n13124;
  reg [63:0] n13126;
  reg [63:0] n13128;
  reg [63:0] n13130;
  reg [4:0] n13131;
  reg n13134;
  wire [31:0] n13135;
  wire n13137;
  wire [31:0] n13138;
  wire [31:0] n13140;
  wire [30:0] n13141;
  wire [63:0] n13142;
  wire [31:0] n13143;
  wire [31:0] n13145;
  wire [30:0] n13146;
  wire [63:0] n13147;
  wire [31:0] n13148;
  wire [31:0] n13150;
  wire [3:0] n13151;
  wire n13157;
  wire n13159;
  wire [63:0] n13160;
  wire [63:0] n13161;
  wire [63:0] n13162;
  wire [63:0] n13163;
  wire [63:0] n13164;
  wire [63:0] n13165;
  wire [63:0] n13166;
  wire [63:0] n13167;
  wire [63:0] n13168;
  wire n13170;
  wire [63:0] n13171;
  wire [63:0] n13172;
  wire [63:0] n13173;
  wire [63:0] n13174;
  wire [63:0] n13175;
  wire [63:0] n13176;
  wire [63:0] n13177;
  wire [63:0] n13178;
  wire [63:0] n13179;
  wire [63:0] n13180;
  wire [63:0] n13181;
  wire [63:0] n13182;
  wire [31:0] n13183;
  wire [31:0] n13185;
  wire [4:0] n13186;
  wire [63:0] n13187;
  wire n13189;
  wire [63:0] n13190;
  wire n13192;
  wire n13193;
  wire [63:0] n13194;
  wire n13196;
  wire [2:0] n13197;
  reg n13201;
  reg [14:0] n13205;
  reg [63:0] n13206;
  wire [2:0] n13208;
  wire [63:0] n13209;
  wire [63:0] n13210;
  wire [63:0] n13211;
  wire [4:0] n13212;
  wire n13213;
  wire [14:0] n13214;
  wire [63:0] n13215;
  wire [63:0] n13216;
  wire [63:0] n13217;
  wire [63:0] n13218;
  wire [2:0] n13219;
  wire [63:0] n13220;
  wire [63:0] n13221;
  wire [63:0] n13222;
  wire [4:0] n13223;
  wire n13224;
  wire n13225;
  wire [14:0] n13226;
  wire [63:0] n13227;
  wire [63:0] n13228;
  wire [63:0] n13229;
  wire [63:0] n13230;
  wire n13232;
  wire n13234;
  wire n13236;
  wire n13237;
  wire n13238;
  wire n13239;
  wire n13240;
  wire [62:0] n13241;
  wire [63:0] n13243;
  wire n13244;
  wire [61:0] n13245;
  wire [63:0] n13247;
  wire [59:0] n13248;
  wire [63:0] n13250;
  wire [14:0] n13253;
  wire [63:0] n13254;
  wire [14:0] n13256;
  wire [63:0] n13257;
  wire [14:0] n13258;
  wire [63:0] n13259;
  wire n13261;
  wire n13262;
  wire [62:0] n13263;
  wire n13265;
  wire n13266;
  wire n13268;
  wire n13269;
  wire n13271;
  wire n13273;
  wire n13274;
  wire n13275;
  wire n13276;
  wire n13278;
  wire n13279;
  wire n13281;
  wire n13282;
  wire n13283;
  wire n13284;
  wire n13285;
  wire n13286;
  wire [1:0] n13287;
  wire [61:0] n13288;
  wire [61:0] n13289;
  wire [61:0] n13290;
  wire [1:0] n13291;
  wire [1:0] n13292;
  wire n13294;
  wire [15:0] n13295;
  wire [79:0] n13296;
  wire n13298;
  wire [7:0] n13299;
  reg [79:0] n13301;
  reg n13305;
  reg n13308;
  reg n13312;
  reg [2:0] n13317;
  reg [63:0] n13319;
  reg [63:0] n13321;
  reg [63:0] n13323;
  reg [4:0] n13325;
  reg n13327;
  reg n13329;
  reg [14:0] n13331;
  wire [61:0] n13332;
  wire [61:0] n13333;
  wire [61:0] n13334;
  wire [61:0] n13335;
  wire [61:0] n13336;
  reg [61:0] n13338;
  wire [1:0] n13339;
  wire [1:0] n13340;
  wire [1:0] n13341;
  wire [1:0] n13342;
  wire [1:0] n13343;
  reg [1:0] n13345;
  reg [79:0] n13349;
  reg [79:0] n13351;
  reg [3:0] n13353;
  reg n13356;
  reg n13359;
  reg n13362;
  reg n13365;
  reg [79:0] n13369;
  reg [79:0] n13371;
  reg [127:0] n13373;
  reg [127:0] n13375;
  reg [127:0] n13377;
  reg [63:0] n13379;
  reg [63:0] n13381;
  reg [63:0] n13383;
  reg [63:0] n13385;
  reg [63:0] n13387;
  reg [63:0] n13389;
  reg [63:0] n13391;
  reg [63:0] n13393;
  reg [63:0] n13395;
  wire [63:0] n13408;
  wire [2:0] n13515;
  reg [2:0] n13516;
  wire n13517;
  wire n13518;
  wire [63:0] n13519;
  reg [63:0] n13520;
  wire n13521;
  wire n13522;
  wire [63:0] n13523;
  reg [63:0] n13524;
  wire n13525;
  wire n13526;
  wire [63:0] n13527;
  reg [63:0] n13528;
  wire n13529;
  wire n13530;
  wire [4:0] n13531;
  reg [4:0] n13532;
  wire n13533;
  wire n13534;
  wire n13535;
  reg n13536;
  wire n13537;
  wire n13538;
  wire n13539;
  reg n13540;
  wire n13541;
  wire n13542;
  wire [14:0] n13543;
  reg [14:0] n13544;
  wire n13545;
  wire n13546;
  wire [63:0] n13547;
  reg [63:0] n13548;
  wire n13553;
  wire n13554;
  wire [79:0] n13555;
  reg [79:0] n13556;
  wire n13557;
  wire n13558;
  wire [79:0] n13559;
  reg [79:0] n13560;
  wire n13561;
  wire n13562;
  wire [3:0] n13563;
  reg [3:0] n13564;
  wire n13565;
  reg n13566;
  wire n13567;
  reg n13568;
  wire n13569;
  reg n13570;
  wire n13571;
  reg n13572;
  wire n13577;
  wire n13578;
  wire [79:0] n13579;
  reg [79:0] n13580;
  wire n13581;
  wire n13582;
  wire [79:0] n13583;
  reg [79:0] n13584;
  wire n13586;
  wire n13587;
  wire [127:0] n13588;
  reg [127:0] n13589;
  wire n13590;
  wire n13591;
  wire [127:0] n13592;
  reg [127:0] n13593;
  wire n13594;
  wire n13595;
  wire [127:0] n13596;
  reg [127:0] n13597;
  wire n13598;
  wire n13599;
  wire [63:0] n13600;
  reg [63:0] n13601;
  wire n13602;
  wire n13603;
  wire [63:0] n13604;
  reg [63:0] n13605;
  wire n13606;
  wire n13607;
  wire [63:0] n13608;
  reg [63:0] n13609;
  wire n13610;
  wire n13611;
  wire [63:0] n13612;
  reg [63:0] n13613;
  wire n13614;
  wire n13615;
  wire [63:0] n13616;
  reg [63:0] n13617;
  wire n13619;
  wire n13620;
  wire [63:0] n13621;
  reg [63:0] n13622;
  wire n13623;
  wire n13624;
  wire [63:0] n13625;
  reg [63:0] n13626;
  wire n13627;
  wire n13628;
  wire [63:0] n13629;
  reg [63:0] n13630;
  wire n13631;
  wire n13632;
  wire [63:0] n13633;
  reg [63:0] n13634;
  wire [79:0] n13635;
  reg [79:0] n13636;
  wire n13637;
  reg n13638;
  wire n13639;
  reg n13640;
  wire n13641;
  reg n13642;
  wire [63:0] n13645; // mem_rd
  assign result = n13636; //(module output)
  assign result_valid = n13638; //(module output)
  assign overflow = trans_overflow; //(module output)
  assign underflow = trans_underflow; //(module output)
  assign inexact = trans_inexact; //(module output)
  assign invalid = trans_invalid; //(module output)
  assign operation_busy = n13640; //(module output)
  assign operation_done = n13642; //(module output)
  /* TG68K_FPU_Transcendental.vhd:102:16  */
  always @*
    trans_state = n13516; // (isignal)
  initial
    trans_state = 3'b000;
  /* TG68K_FPU_Transcendental.vhd:126:16  */
  assign cordic_x = n13520; // (signal)
  /* TG68K_FPU_Transcendental.vhd:126:26  */
  assign cordic_y = n13524; // (signal)
  /* TG68K_FPU_Transcendental.vhd:126:36  */
  assign cordic_z = n13528; // (signal)
  /* TG68K_FPU_Transcendental.vhd:127:16  */
  assign cordic_iteration = n13532; // (signal)
  /* TG68K_FPU_Transcendental.vhd:128:16  */
  assign cordic_mode = n13536; // (signal)
  /* TG68K_FPU_Transcendental.vhd:131:16  */
  assign input_sign = n11071; // (signal)
  /* TG68K_FPU_Transcendental.vhd:132:16  */
  assign input_exp = n11072; // (signal)
  /* TG68K_FPU_Transcendental.vhd:133:16  */
  assign input_mant = n11073; // (signal)
  /* TG68K_FPU_Transcendental.vhd:134:16  */
  assign input_zero = n11083; // (signal)
  /* TG68K_FPU_Transcendental.vhd:135:16  */
  assign input_inf = n11095; // (signal)
  /* TG68K_FPU_Transcendental.vhd:136:16  */
  assign input_nan = n11108; // (signal)
  /* TG68K_FPU_Transcendental.vhd:139:16  */
  assign result_sign = n13540; // (signal)
  /* TG68K_FPU_Transcendental.vhd:140:16  */
  assign result_exp = n13544; // (signal)
  /* TG68K_FPU_Transcendental.vhd:141:16  */
  assign result_mant = n13548; // (signal)
  /* TG68K_FPU_Transcendental.vhd:145:16  */
  assign series_term = n13556; // (signal)
  /* TG68K_FPU_Transcendental.vhd:146:16  */
  assign series_sum = n13560; // (signal)
  /* TG68K_FPU_Transcendental.vhd:147:16  */
  assign iteration_count = n13564; // (signal)
  /* TG68K_FPU_Transcendental.vhd:150:16  */
  assign trans_overflow = n13566; // (signal)
  /* TG68K_FPU_Transcendental.vhd:151:16  */
  assign trans_underflow = n13568; // (signal)
  /* TG68K_FPU_Transcendental.vhd:152:16  */
  assign trans_inexact = n13570; // (signal)
  /* TG68K_FPU_Transcendental.vhd:153:16  */
  assign trans_invalid = n13572; // (signal)
  /* TG68K_FPU_Transcendental.vhd:157:16  */
  assign exp_argument = n13580; // (signal)
  /* TG68K_FPU_Transcendental.vhd:158:16  */
  assign log_argument = n13584; // (signal)
  /* TG68K_FPU_Transcendental.vhd:162:16  */
  assign x_squared = n13589; // (signal)
  /* TG68K_FPU_Transcendental.vhd:163:16  */
  assign x_cubed = n13593; // (signal)
  /* TG68K_FPU_Transcendental.vhd:164:16  */
  assign x_fifth = n13597; // (signal)
  /* TG68K_FPU_Transcendental.vhd:165:16  */
  assign x3_div6 = n13601; // (signal)
  /* TG68K_FPU_Transcendental.vhd:168:16  */
  assign cordic_shift_x = n13605; // (signal)
  /* TG68K_FPU_Transcendental.vhd:169:16  */
  assign cordic_shift_y = n13609; // (signal)
  /* TG68K_FPU_Transcendental.vhd:170:16  */
  assign cordic_atan_val = n13613; // (signal)
  /* TG68K_FPU_Transcendental.vhd:171:16  */
  assign x5_div120 = n13617; // (signal)
  /* TG68K_FPU_Transcendental.vhd:175:16  */
  assign x_n = n13622; // (signal)
  /* TG68K_FPU_Transcendental.vhd:176:16  */
  assign a_div_x_n = n13626; // (signal)
  /* TG68K_FPU_Transcendental.vhd:177:16  */
  assign x_next = n13630; // (signal)
  /* TG68K_FPU_Transcendental.vhd:178:16  */
  assign final_mant = n13634; // (signal)
  /* TG68K_FPU_Transcendental.vhd:185:38  */
  assign n11071 = operand[79]; // extract
  /* TG68K_FPU_Transcendental.vhd:186:37  */
  assign n11072 = operand[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:187:38  */
  assign n11073 = operand[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:190:27  */
  assign n11074 = operand[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:190:42  */
  assign n11076 = n11074 == 15'b000000000000000;
  /* TG68K_FPU_Transcendental.vhd:190:73  */
  assign n11077 = operand[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:190:87  */
  assign n11079 = n11077 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:190:62  */
  assign n11080 = n11079 & n11076;
  /* TG68K_FPU_Transcendental.vhd:190:17  */
  assign n11083 = n11080 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:196:27  */
  assign n11084 = operand[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:196:42  */
  assign n11086 = n11084 == 15'b111111111111111;
  /* TG68K_FPU_Transcendental.vhd:196:73  */
  assign n11087 = operand[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:196:62  */
  assign n11088 = n11087 & n11086;
  /* TG68K_FPU_Transcendental.vhd:196:95  */
  assign n11089 = operand[62:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:196:109  */
  assign n11091 = n11089 == 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:196:84  */
  assign n11092 = n11091 & n11088;
  /* TG68K_FPU_Transcendental.vhd:196:17  */
  assign n11095 = n11092 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:202:27  */
  assign n11096 = operand[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:202:42  */
  assign n11098 = n11096 == 15'b111111111111111;
  /* TG68K_FPU_Transcendental.vhd:202:78  */
  assign n11099 = operand[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:202:100  */
  assign n11100 = operand[62:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:202:114  */
  assign n11102 = n11100 == 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:202:89  */
  assign n11103 = n11102 & n11099;
  /* TG68K_FPU_Transcendental.vhd:202:66  */
  assign n11104 = ~n11103;
  /* TG68K_FPU_Transcendental.vhd:202:62  */
  assign n11105 = n11104 & n11098;
  /* TG68K_FPU_Transcendental.vhd:202:17  */
  assign n11108 = n11105 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:219:27  */
  assign n11111 = ~nreset;
  /* TG68K_FPU_Transcendental.vhd:242:49  */
  assign n11115 = start_operation ? 1'b1 : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:242:49  */
  assign n11118 = start_operation ? 3'b001 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:242:49  */
  assign n11122 = start_operation ? 4'b0000 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:233:41  */
  assign n11124 = trans_state == 3'b000;
  /* TG68K_FPU_Transcendental.vhd:260:65  */
  assign n11126 = operation_code == 7'b0001110;
  /* TG68K_FPU_Transcendental.vhd:260:78  */
  assign n11128 = operation_code == 7'b0011101;
  /* TG68K_FPU_Transcendental.vhd:260:78  */
  assign n11129 = n11126 | n11128;
  /* TG68K_FPU_Transcendental.vhd:260:88  */
  assign n11131 = operation_code == 7'b0001111;
  /* TG68K_FPU_Transcendental.vhd:260:88  */
  assign n11132 = n11129 | n11131;
  /* TG68K_FPU_Transcendental.vhd:267:87  */
  assign n11133 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:267:73  */
  assign n11136 = n11133 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : 64'b1100000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:267:73  */
  assign n11138 = n11133 ? trans_invalid : 1'b1;
  /* TG68K_FPU_Transcendental.vhd:266:65  */
  assign n11140 = operation_code == 7'b0000100;
  assign n11141 = {n11140, n11132};
  /* TG68K_FPU_Transcendental.vhd:259:57  */
  always @*
    case (n11141)
      2'b10: n11144 = 1'b0;
      2'b01: n11144 = 1'b0;
      default: n11144 = input_sign;
    endcase
  /* TG68K_FPU_Transcendental.vhd:259:57  */
  always @*
    case (n11141)
      2'b10: n11147 = 15'b111111111111111;
      2'b01: n11147 = 15'b111111111111111;
      default: n11147 = input_exp;
    endcase
  /* TG68K_FPU_Transcendental.vhd:259:57  */
  always @*
    case (n11141)
      2'b10: n11149 = n11136;
      2'b01: n11149 = 64'b1100000000000000000000000000000000000000000000000000000000000000;
      default: n11149 = input_mant;
    endcase
  /* TG68K_FPU_Transcendental.vhd:259:57  */
  always @*
    case (n11141)
      2'b10: n11151 = n11138;
      2'b01: n11151 = 1'b1;
      default: n11151 = trans_invalid;
    endcase
  /* TG68K_FPU_Transcendental.vhd:257:49  */
  assign n11154 = input_inf ? 3'b111 : 3'b010;
  /* TG68K_FPU_Transcendental.vhd:257:49  */
  assign n11155 = input_inf ? n11144 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:257:49  */
  assign n11156 = input_inf ? n11147 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:257:49  */
  assign n11157 = input_inf ? n11149 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:257:49  */
  assign n11158 = input_inf ? n11151 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:251:49  */
  assign n11160 = input_nan ? 3'b111 : n11154;
  /* TG68K_FPU_Transcendental.vhd:251:49  */
  assign n11161 = input_nan ? input_sign : n11155;
  /* TG68K_FPU_Transcendental.vhd:251:49  */
  assign n11163 = input_nan ? 15'b111111111111111 : n11156;
  /* TG68K_FPU_Transcendental.vhd:251:49  */
  assign n11164 = input_nan ? input_mant : n11157;
  /* TG68K_FPU_Transcendental.vhd:251:49  */
  assign n11165 = input_nan ? trans_invalid : n11158;
  /* TG68K_FPU_Transcendental.vhd:249:41  */
  assign n11167 = trans_state == 3'b001;
  /* TG68K_FPU_Transcendental.vhd:294:100  */
  assign n11168 = ~input_zero;
  /* TG68K_FPU_Transcendental.vhd:294:85  */
  assign n11169 = n11168 & input_sign;
  /* TG68K_FPU_Transcendental.vhd:301:65  */
  assign n11172 = input_zero ? 3'b111 : 3'b011;
  /* TG68K_FPU_Transcendental.vhd:301:65  */
  assign n11173 = input_zero ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:301:65  */
  assign n11175 = input_zero ? 15'b000000000000000 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:301:65  */
  assign n11177 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:294:65  */
  assign n11179 = n11169 ? 3'b111 : n11172;
  /* TG68K_FPU_Transcendental.vhd:294:65  */
  assign n11181 = n11169 ? 1'b0 : n11173;
  /* TG68K_FPU_Transcendental.vhd:294:65  */
  assign n11183 = n11169 ? 15'b111111111111111 : n11175;
  /* TG68K_FPU_Transcendental.vhd:294:65  */
  assign n11185 = n11169 ? 64'b1100000000000000000000000000000000000000000000000000000000000000 : n11177;
  /* TG68K_FPU_Transcendental.vhd:294:65  */
  assign n11187 = n11169 ? 1'b1 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:293:57  */
  assign n11189 = operation_code == 7'b0000100;
  /* TG68K_FPU_Transcendental.vhd:314:91  */
  assign n11191 = operation_code == 7'b0001110;
  /* TG68K_FPU_Transcendental.vhd:314:119  */
  assign n11193 = operation_code == 7'b0001111;
  /* TG68K_FPU_Transcendental.vhd:314:101  */
  assign n11194 = n11191 | n11193;
  /* TG68K_FPU_Transcendental.vhd:314:73  */
  assign n11196 = n11194 ? input_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:314:73  */
  assign n11199 = n11194 ? 15'b000000000000000 : 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:314:73  */
  assign n11202 = n11194 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:312:65  */
  assign n11205 = input_zero ? 3'b111 : 3'b011;
  /* TG68K_FPU_Transcendental.vhd:312:65  */
  assign n11206 = input_zero ? n11196 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:312:65  */
  assign n11207 = input_zero ? n11199 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:312:65  */
  assign n11208 = input_zero ? n11202 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:311:57  */
  assign n11211 = operation_code == 7'b0001110;
  /* TG68K_FPU_Transcendental.vhd:311:70  */
  assign n11213 = operation_code == 7'b0011101;
  /* TG68K_FPU_Transcendental.vhd:311:70  */
  assign n11214 = n11211 | n11213;
  /* TG68K_FPU_Transcendental.vhd:311:80  */
  assign n11216 = operation_code == 7'b0001111;
  /* TG68K_FPU_Transcendental.vhd:311:80  */
  assign n11217 = n11214 | n11216;
  /* TG68K_FPU_Transcendental.vhd:338:65  */
  assign n11220 = input_zero ? 3'b111 : 3'b011;
  /* TG68K_FPU_Transcendental.vhd:338:65  */
  assign n11222 = input_zero ? 1'b1 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:338:65  */
  assign n11224 = input_zero ? 15'b111111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:338:65  */
  assign n11226 = input_zero ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:338:65  */
  assign n11227 = input_zero ? log_argument : operand;
  /* TG68K_FPU_Transcendental.vhd:331:65  */
  assign n11229 = input_sign ? 3'b111 : n11220;
  /* TG68K_FPU_Transcendental.vhd:331:65  */
  assign n11231 = input_sign ? 1'b0 : n11222;
  /* TG68K_FPU_Transcendental.vhd:331:65  */
  assign n11233 = input_sign ? 15'b111111111111111 : n11224;
  /* TG68K_FPU_Transcendental.vhd:331:65  */
  assign n11235 = input_sign ? 64'b1100000000000000000000000000000000000000000000000000000000000000 : n11226;
  /* TG68K_FPU_Transcendental.vhd:331:65  */
  assign n11237 = input_sign ? 1'b1 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:331:65  */
  assign n11238 = input_sign ? log_argument : n11227;
  /* TG68K_FPU_Transcendental.vhd:330:57  */
  assign n11240 = operation_code == 7'b0010100;
  /* TG68K_FPU_Transcendental.vhd:330:71  */
  assign n11242 = operation_code == 7'b0010110;
  /* TG68K_FPU_Transcendental.vhd:330:71  */
  assign n11243 = n11240 | n11242;
  /* TG68K_FPU_Transcendental.vhd:330:82  */
  assign n11245 = operation_code == 7'b0010101;
  /* TG68K_FPU_Transcendental.vhd:330:82  */
  assign n11246 = n11243 | n11245;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n11247 = {n11246, n11217, n11189};
  /* TG68K_FPU_Transcendental.vhd:292:49  */
  always @*
    case (n11247)
      3'b100: n11249 = n11229;
      3'b010: n11249 = n11205;
      3'b001: n11249 = n11179;
      default: n11249 = 3'b011;
    endcase
  /* TG68K_FPU_Transcendental.vhd:292:49  */
  always @*
    case (n11247)
      3'b100: n11250 = n11231;
      3'b010: n11250 = n11206;
      3'b001: n11250 = n11181;
      default: n11250 = result_sign;
    endcase
  /* TG68K_FPU_Transcendental.vhd:292:49  */
  always @*
    case (n11247)
      3'b100: n11251 = n11233;
      3'b010: n11251 = n11207;
      3'b001: n11251 = n11183;
      default: n11251 = result_exp;
    endcase
  /* TG68K_FPU_Transcendental.vhd:292:49  */
  always @*
    case (n11247)
      3'b100: n11252 = n11235;
      3'b010: n11252 = n11208;
      3'b001: n11252 = n11185;
      default: n11252 = result_mant;
    endcase
  /* TG68K_FPU_Transcendental.vhd:292:49  */
  always @*
    case (n11247)
      3'b100: n11253 = n11237;
      3'b010: n11253 = trans_invalid;
      3'b001: n11253 = n11187;
      default: n11253 = trans_invalid;
    endcase
  /* TG68K_FPU_Transcendental.vhd:292:49  */
  always @*
    case (n11247)
      3'b100: n11255 = n11238;
      3'b010: n11255 = log_argument;
      3'b001: n11255 = log_argument;
      default: n11255 = log_argument;
    endcase
  /* TG68K_FPU_Transcendental.vhd:290:41  */
  assign n11257 = trans_state == 3'b010;
  /* TG68K_FPU_Transcendental.vhd:359:84  */
  assign n11258 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:359:84  */
  assign n11260 = n11258 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:362:85  */
  assign n11261 = input_exp[0]; // extract
  /* TG68K_FPU_Transcendental.vhd:362:89  */
  assign n11262 = ~n11261;
  /* TG68K_FPU_Transcendental.vhd:364:144  */
  assign n11264 = input_exp - 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:364:112  */
  assign n11266 = n11264 >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:364:156  */
  assign n11268 = n11266 + 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:367:144  */
  assign n11270 = input_exp - 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:367:152  */
  assign n11272 = n11270 + 15'b000000000000001;
  /* TG68K_FPU_Transcendental.vhd:367:112  */
  assign n11274 = n11272 >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:367:160  */
  assign n11276 = n11274 + 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:362:73  */
  assign n11277 = n11262 ? n11268 : n11276;
  /* TG68K_FPU_Transcendental.vhd:371:108  */
  assign n11278 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:371:108  */
  assign n11280 = n11278 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:371:92  */
  assign n11281 = n11280[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:372:87  */
  assign n11282 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:372:87  */
  assign n11284 = $signed(n11282) < $signed(32'b00000000000000000000000000001000);
  /* TG68K_FPU_Transcendental.vhd:375:88  */
  assign n11285 = x_n[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:375:104  */
  assign n11287 = $unsigned(n11285) > $unsigned(16'b0000000000000000);
  /* TG68K_FPU_Transcendental.vhd:378:115  */
  assign n11288 = input_mant[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:378:131  */
  assign n11289 = {16'b0, n11288};  //  uext
  /* TG68K_FPU_Transcendental.vhd:378:131  */
  assign n11291 = $signed(n11289) * $signed(32'b00000000000000010000000000000000); // smul
  /* TG68K_FPU_Transcendental.vhd:378:153  */
  assign n11292 = x_n[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:378:139  */
  assign n11293 = {16'b0, n11292};  //  uext
  /* TG68K_FPU_Transcendental.vhd:378:139  */
  assign n11294 = n11291 / n11293; // udiv
  /* TG68K_FPU_Transcendental.vhd:378:89  */
  assign n11295 = {32'b0, n11294};  //  uext
  /* TG68K_FPU_Transcendental.vhd:375:73  */
  assign n11296 = n11287 ? n11295 : input_mant;
  /* TG68K_FPU_Transcendental.vhd:385:126  */
  assign n11297 = x_n + a_div_x_n;
  /* TG68K_FPU_Transcendental.vhd:385:100  */
  assign n11299 = n11297 >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:387:108  */
  assign n11300 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:387:108  */
  assign n11302 = n11300 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:387:92  */
  assign n11303 = n11302[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:394:85  */
  assign n11304 = input_exp[0]; // extract
  /* TG68K_FPU_Transcendental.vhd:399:89  */
  assign n11306 = x_n >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:398:103  */
  assign n11307 = x_n + n11306;
  /* TG68K_FPU_Transcendental.vhd:400:89  */
  assign n11309 = x_n >> 31'b0000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:399:119  */
  assign n11310 = n11307 + n11309;
  /* TG68K_FPU_Transcendental.vhd:401:89  */
  assign n11312 = x_n >> 31'b0000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:400:119  */
  assign n11313 = n11310 - n11312;
  /* TG68K_FPU_Transcendental.vhd:394:73  */
  assign n11314 = n11304 ? n11313 : x_n;
  /* TG68K_FPU_Transcendental.vhd:409:86  */
  assign n11315 = final_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:409:91  */
  assign n11316 = ~n11315;
  /* TG68K_FPU_Transcendental.vhd:411:106  */
  assign n11317 = final_mant[62:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:411:120  */
  assign n11319 = {n11317, 1'b0};
  /* TG68K_FPU_Transcendental.vhd:412:133  */
  assign n11321 = result_exp - 15'b000000000000001;
  /* TG68K_FPU_Transcendental.vhd:409:73  */
  assign n11322 = n11316 ? n11321 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:409:73  */
  assign n11323 = n11316 ? n11319 : final_mant;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11325 = n11284 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11327 = n11284 ? result_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11328 = n11284 ? result_exp : n11322;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11329 = n11284 ? result_mant : n11323;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11330 = n11284 ? n11303 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11332 = n11284 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11333 = n11284 ? x_next : x_n;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11334 = n11284 ? n11296 : a_div_x_n;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11335 = n11284 ? n11299 : x_next;
  /* TG68K_FPU_Transcendental.vhd:372:65  */
  assign n11336 = n11284 ? final_mant : n11314;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11337 = n11260 ? trans_state : n11325;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11338 = n11260 ? result_sign : n11327;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11339 = n11260 ? n11277 : n11328;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11340 = n11260 ? result_mant : n11329;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11341 = n11260 ? n11281 : n11330;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11342 = n11260 ? trans_inexact : n11332;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11344 = n11260 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n11333;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11345 = n11260 ? a_div_x_n : n11334;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11346 = n11260 ? x_next : n11335;
  /* TG68K_FPU_Transcendental.vhd:359:65  */
  assign n11347 = n11260 ? final_mant : n11336;
  /* TG68K_FPU_Transcendental.vhd:357:57  */
  assign n11349 = operation_code == 7'b0000100;
  /* TG68K_FPU_Transcendental.vhd:422:88  */
  assign n11351 = $unsigned(input_exp) < $unsigned(15'b011111111110101);
  /* TG68K_FPU_Transcendental.vhd:422:65  */
  assign n11354 = n11351 ? 3'b110 : 3'b101;
  /* TG68K_FPU_Transcendental.vhd:422:65  */
  assign n11356 = n11351 ? cordic_iteration : 5'b00000;
  /* TG68K_FPU_Transcendental.vhd:422:65  */
  assign n11357 = n11351 ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:422:65  */
  assign n11358 = n11351 ? input_exp : result_exp;
  /* TG68K_FPU_Transcendental.vhd:422:65  */
  assign n11359 = n11351 ? input_mant : result_mant;
  /* TG68K_FPU_Transcendental.vhd:420:57  */
  assign n11361 = operation_code == 7'b0001110;
  /* TG68K_FPU_Transcendental.vhd:436:88  */
  assign n11363 = $unsigned(input_exp) < $unsigned(15'b011111111110101);
  /* TG68K_FPU_Transcendental.vhd:436:65  */
  assign n11366 = n11363 ? 3'b110 : 3'b101;
  /* TG68K_FPU_Transcendental.vhd:436:65  */
  assign n11368 = n11363 ? cordic_iteration : 5'b00000;
  /* TG68K_FPU_Transcendental.vhd:436:65  */
  assign n11370 = n11363 ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:436:65  */
  assign n11372 = n11363 ? 15'b011111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:436:65  */
  assign n11374 = n11363 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:434:57  */
  assign n11376 = operation_code == 7'b0011101;
  /* TG68K_FPU_Transcendental.vhd:450:84  */
  assign n11377 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:450:84  */
  assign n11379 = n11377 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:452:96  */
  assign n11381 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:452:135  */
  assign n11382 = input_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:452:121  */
  assign n11383 = n11382 & n11381;
  /* TG68K_FPU_Transcendental.vhd:452:160  */
  assign n11384 = input_mant[62:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:452:174  */
  assign n11386 = n11384 == 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:452:146  */
  assign n11387 = n11386 & n11383;
  /* TG68K_FPU_Transcendental.vhd:460:116  */
  assign n11388 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:460:116  */
  assign n11390 = n11388 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:460:100  */
  assign n11391 = n11390[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:452:73  */
  assign n11393 = n11387 ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:452:73  */
  assign n11395 = n11387 ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:452:73  */
  assign n11397 = n11387 ? 15'b000000000000000 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:452:73  */
  assign n11399 = n11387 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:452:73  */
  assign n11400 = n11387 ? iteration_count : n11391;
  /* TG68K_FPU_Transcendental.vhd:452:73  */
  assign n11401 = n11387 ? log_argument : operand;
  /* TG68K_FPU_Transcendental.vhd:462:87  */
  assign n11402 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:462:87  */
  assign n11404 = $signed(n11402) <= $signed(32'b00000000000000000000000000000110);
  /* TG68K_FPU_Transcendental.vhd:465:92  */
  assign n11405 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:465:92  */
  assign n11407 = n11405 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:467:104  */
  assign n11409 = $unsigned(input_exp) >= $unsigned(15'b011111111111111);
  /* TG68K_FPU_Transcendental.vhd:470:125  */
  assign n11411 = input_exp - 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:470:134  */
  assign n11412 = {16'b0, n11411};  //  uext
  /* TG68K_FPU_Transcendental.vhd:470:134  */
  assign n11415 = n11412 * 31'b0000000000000001011000101110010; // umul
  /* TG68K_FPU_Transcendental.vhd:470:97  */
  assign n11416 = {49'b0, n11415};  //  uext
  /* TG68K_FPU_Transcendental.vhd:475:119  */
  assign n11418 = 15'b011111111111111 - input_exp;
  /* TG68K_FPU_Transcendental.vhd:475:142  */
  assign n11419 = {16'b0, n11418};  //  uext
  /* TG68K_FPU_Transcendental.vhd:475:142  */
  assign n11422 = n11419 * 31'b0000000000000001011000101110010; // umul
  /* TG68K_FPU_Transcendental.vhd:475:104  */
  assign n11423 = -n11422;
  /* TG68K_FPU_Transcendental.vhd:475:97  */
  assign n11424 = {{49{n11423[30]}}, n11423}; // sext
  /* TG68K_FPU_Transcendental.vhd:467:81  */
  assign n11425 = n11409 ? n11416 : n11424;
  /* TG68K_FPU_Transcendental.vhd:478:95  */
  assign n11426 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:478:95  */
  assign n11428 = $signed(n11426) <= $signed(32'b00000000000000000000000000000100);
  /* TG68K_FPU_Transcendental.vhd:482:94  */
  assign n11429 = input_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:484:147  */
  assign n11430 = input_mant[62:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:484:121  */
  assign n11431 = {17'b0, n11430};  //  uext
  /* TG68K_FPU_Transcendental.vhd:486:141  */
  assign n11432 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:478:73  */
  assign n11433 = n11435 ? n11431 : series_term;
  /* TG68K_FPU_Transcendental.vhd:478:73  */
  assign n11434 = n11436 ? n11432 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:478:73  */
  assign n11435 = n11429 & n11428;
  /* TG68K_FPU_Transcendental.vhd:478:73  */
  assign n11436 = n11429 & n11428;
  /* TG68K_FPU_Transcendental.vhd:465:73  */
  assign n11437 = n11407 ? series_term : n11433;
  /* TG68K_FPU_Transcendental.vhd:465:73  */
  assign n11438 = n11407 ? n11425 : n11434;
  /* TG68K_FPU_Transcendental.vhd:492:108  */
  assign n11439 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:492:108  */
  assign n11441 = n11439 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:492:92  */
  assign n11442 = n11441[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:496:95  */
  assign n11443 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:496:111  */
  assign n11445 = n11443 == 15'b000000000000000;
  /* TG68K_FPU_Transcendental.vhd:496:129  */
  assign n11446 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:496:143  */
  assign n11448 = n11446 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:496:115  */
  assign n11449 = n11448 & n11445;
  /* TG68K_FPU_Transcendental.vhd:503:106  */
  assign n11450 = series_sum[79]; // extract
  /* TG68K_FPU_Transcendental.vhd:504:105  */
  assign n11451 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:505:106  */
  assign n11452 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:496:73  */
  assign n11454 = n11449 ? 1'b0 : n11450;
  /* TG68K_FPU_Transcendental.vhd:496:73  */
  assign n11456 = n11449 ? 15'b000000000000000 : n11451;
  /* TG68K_FPU_Transcendental.vhd:496:73  */
  assign n11458 = n11449 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n11452;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11460 = n11404 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11461 = n11404 ? result_sign : n11454;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11462 = n11404 ? result_exp : n11456;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11463 = n11404 ? result_mant : n11458;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11464 = n11404 ? n11437 : series_term;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11465 = n11404 ? n11438 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11466 = n11404 ? n11442 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:462:65  */
  assign n11468 = n11404 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11469 = n11379 ? n11393 : n11460;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11470 = n11379 ? n11395 : n11461;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11471 = n11379 ? n11397 : n11462;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11472 = n11379 ? n11399 : n11463;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11473 = n11379 ? series_term : n11464;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11474 = n11379 ? series_sum : n11465;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11475 = n11379 ? n11400 : n11466;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11476 = n11379 ? trans_inexact : n11468;
  /* TG68K_FPU_Transcendental.vhd:450:65  */
  assign n11477 = n11379 ? n11401 : log_argument;
  /* TG68K_FPU_Transcendental.vhd:448:57  */
  assign n11479 = operation_code == 7'b0010100;
  /* TG68K_FPU_Transcendental.vhd:512:84  */
  assign n11480 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:512:84  */
  assign n11482 = $signed(n11480) < $signed(32'b00000000000000000000000000000110);
  /* TG68K_FPU_Transcendental.vhd:513:108  */
  assign n11483 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:513:108  */
  assign n11485 = n11483 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:513:92  */
  assign n11486 = n11485[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:517:96  */
  assign n11488 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:517:135  */
  assign n11489 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:517:150  */
  assign n11491 = n11489 == 32'b10000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:517:121  */
  assign n11492 = n11491 & n11488;
  /* TG68K_FPU_Transcendental.vhd:526:140  */
  assign n11494 = input_exp - 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:526:113  */
  assign n11495 = {49'b0, n11494};  //  uext
  /* TG68K_FPU_Transcendental.vhd:517:73  */
  assign n11498 = n11492 ? 15'b000000000000000 : 15'b011111111111101;
  /* TG68K_FPU_Transcendental.vhd:517:73  */
  assign n11500 = n11492 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n11495;
  /* TG68K_FPU_Transcendental.vhd:512:65  */
  assign n11502 = n11482 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:512:65  */
  assign n11504 = n11482 ? result_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:512:65  */
  assign n11505 = n11482 ? result_exp : n11498;
  /* TG68K_FPU_Transcendental.vhd:512:65  */
  assign n11506 = n11482 ? result_mant : n11500;
  /* TG68K_FPU_Transcendental.vhd:512:65  */
  assign n11507 = n11482 ? n11486 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:510:57  */
  assign n11509 = operation_code == 7'b0010101;
  /* TG68K_FPU_Transcendental.vhd:534:84  */
  assign n11510 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:534:84  */
  assign n11512 = $signed(n11510) < $signed(32'b00000000000000000000000000000110);
  /* TG68K_FPU_Transcendental.vhd:535:108  */
  assign n11513 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:535:108  */
  assign n11515 = n11513 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:535:92  */
  assign n11516 = n11515[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:539:96  */
  assign n11518 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:539:135  */
  assign n11519 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:539:150  */
  assign n11521 = n11519 == 32'b10000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:539:121  */
  assign n11522 = n11521 & n11518;
  /* TG68K_FPU_Transcendental.vhd:548:140  */
  assign n11524 = input_exp - 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:548:113  */
  assign n11525 = {49'b0, n11524};  //  uext
  /* TG68K_FPU_Transcendental.vhd:539:73  */
  assign n11528 = n11522 ? 15'b000000000000000 : 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:539:73  */
  assign n11530 = n11522 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n11525;
  /* TG68K_FPU_Transcendental.vhd:534:65  */
  assign n11532 = n11512 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:534:65  */
  assign n11534 = n11512 ? result_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:534:65  */
  assign n11535 = n11512 ? result_exp : n11528;
  /* TG68K_FPU_Transcendental.vhd:534:65  */
  assign n11536 = n11512 ? result_mant : n11530;
  /* TG68K_FPU_Transcendental.vhd:534:65  */
  assign n11537 = n11512 ? n11516 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:532:57  */
  assign n11539 = operation_code == 7'b0010110;
  /* TG68K_FPU_Transcendental.vhd:557:84  */
  assign n11540 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:557:84  */
  assign n11542 = n11540 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:568:116  */
  assign n11543 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:568:116  */
  assign n11545 = n11543 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:568:100  */
  assign n11546 = n11545[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:559:73  */
  assign n11548 = input_zero ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:559:73  */
  assign n11549 = input_zero ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:559:73  */
  assign n11551 = input_zero ? 15'b000000000000000 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:559:73  */
  assign n11553 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:559:73  */
  assign n11554 = input_zero ? series_sum : operand;
  /* TG68K_FPU_Transcendental.vhd:559:73  */
  assign n11555 = input_zero ? iteration_count : n11546;
  /* TG68K_FPU_Transcendental.vhd:570:87  */
  assign n11556 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:570:87  */
  assign n11558 = $signed(n11556) <= $signed(32'b00000000000000000000000000001000);
  /* TG68K_FPU_Transcendental.vhd:572:92  */
  assign n11559 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:572:92  */
  assign n11561 = n11559 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:575:115  */
  assign n11562 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:575:152  */
  assign n11563 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:575:131  */
  assign n11564 = {32'b0, n11562};  //  uext
  /* TG68K_FPU_Transcendental.vhd:575:131  */
  assign n11565 = {32'b0, n11563};  //  uext
  /* TG68K_FPU_Transcendental.vhd:575:131  */
  assign n11566 = n11564 * n11565; // umul
  /* TG68K_FPU_Transcendental.vhd:575:89  */
  assign n11567 = {64'b0, n11566};  //  uext
  /* TG68K_FPU_Transcendental.vhd:577:95  */
  assign n11568 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:577:95  */
  assign n11570 = n11568 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:580:114  */
  assign n11571 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:580:152  */
  assign n11572 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:580:131  */
  assign n11573 = {32'b0, n11571};  //  uext
  /* TG68K_FPU_Transcendental.vhd:580:131  */
  assign n11574 = {32'b0, n11572};  //  uext
  /* TG68K_FPU_Transcendental.vhd:580:131  */
  assign n11575 = n11573 * n11574; // umul
  /* TG68K_FPU_Transcendental.vhd:580:89  */
  assign n11576 = {64'b0, n11575};  //  uext
  /* TG68K_FPU_Transcendental.vhd:582:95  */
  assign n11577 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:582:95  */
  assign n11579 = n11577 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:584:132  */
  assign n11580 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:584:149  */
  assign n11582 = n11580 / 32'b00000000000000000000000000000011; // udiv
  /* TG68K_FPU_Transcendental.vhd:584:109  */
  assign n11583 = {32'b0, n11582};  //  uext
  /* TG68K_FPU_Transcendental.vhd:585:95  */
  assign n11584 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:585:95  */
  assign n11586 = n11584 == 32'b00000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:588:89  */
  assign n11587 = {16'b0, x3_div6};  //  uext
  /* TG68K_FPU_Transcendental.vhd:587:133  */
  assign n11588 = series_sum + n11587;
  /* TG68K_FPU_Transcendental.vhd:589:95  */
  assign n11589 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:589:95  */
  assign n11591 = n11589 == 32'b00000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:592:112  */
  assign n11592 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:592:149  */
  assign n11593 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:592:129  */
  assign n11594 = {32'b0, n11592};  //  uext
  /* TG68K_FPU_Transcendental.vhd:592:129  */
  assign n11595 = {32'b0, n11593};  //  uext
  /* TG68K_FPU_Transcendental.vhd:592:129  */
  assign n11596 = n11594 * n11595; // umul
  /* TG68K_FPU_Transcendental.vhd:592:89  */
  assign n11597 = {64'b0, n11596};  //  uext
  /* TG68K_FPU_Transcendental.vhd:594:95  */
  assign n11598 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:594:95  */
  assign n11600 = n11598 == 32'b00000000000000000000000000000110;
  /* TG68K_FPU_Transcendental.vhd:596:146  */
  assign n11601 = x_fifth[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:596:163  */
  assign n11602 = {64'b0, n11601};  //  uext
  /* TG68K_FPU_Transcendental.vhd:596:163  */
  assign n11604 = $signed(n11602) * $signed(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010); // smul
  /* TG68K_FPU_Transcendental.vhd:596:118  */
  assign n11606 = n11604 >> 31'b0000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:596:111  */
  assign n11607 = n11606[63:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:597:95  */
  assign n11608 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:597:95  */
  assign n11610 = n11608 == 32'b00000000000000000000000000000111;
  /* TG68K_FPU_Transcendental.vhd:600:89  */
  assign n11611 = {16'b0, x5_div120};  //  uext
  /* TG68K_FPU_Transcendental.vhd:599:133  */
  assign n11612 = series_sum + n11611;
  /* TG68K_FPU_Transcendental.vhd:597:73  */
  assign n11613 = n11610 ? n11612 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:594:73  */
  assign n11614 = n11600 ? series_sum : n11613;
  /* TG68K_FPU_Transcendental.vhd:594:73  */
  assign n11615 = n11600 ? n11607 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:589:73  */
  assign n11616 = n11591 ? series_sum : n11614;
  /* TG68K_FPU_Transcendental.vhd:589:73  */
  assign n11617 = n11591 ? n11597 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:589:73  */
  assign n11618 = n11591 ? x5_div120 : n11615;
  /* TG68K_FPU_Transcendental.vhd:585:73  */
  assign n11619 = n11586 ? n11588 : n11616;
  /* TG68K_FPU_Transcendental.vhd:585:73  */
  assign n11620 = n11586 ? x_fifth : n11617;
  /* TG68K_FPU_Transcendental.vhd:585:73  */
  assign n11621 = n11586 ? x5_div120 : n11618;
  /* TG68K_FPU_Transcendental.vhd:582:73  */
  assign n11622 = n11579 ? series_sum : n11619;
  /* TG68K_FPU_Transcendental.vhd:582:73  */
  assign n11623 = n11579 ? x_fifth : n11620;
  /* TG68K_FPU_Transcendental.vhd:582:73  */
  assign n11624 = n11579 ? n11583 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:582:73  */
  assign n11625 = n11579 ? x5_div120 : n11621;
  /* TG68K_FPU_Transcendental.vhd:577:73  */
  assign n11626 = n11570 ? series_sum : n11622;
  /* TG68K_FPU_Transcendental.vhd:577:73  */
  assign n11627 = n11570 ? n11576 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:577:73  */
  assign n11628 = n11570 ? x_fifth : n11623;
  /* TG68K_FPU_Transcendental.vhd:577:73  */
  assign n11629 = n11570 ? x3_div6 : n11624;
  /* TG68K_FPU_Transcendental.vhd:577:73  */
  assign n11630 = n11570 ? x5_div120 : n11625;
  /* TG68K_FPU_Transcendental.vhd:572:73  */
  assign n11631 = n11561 ? series_sum : n11626;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11632 = n11659 ? n11567 : x_squared;
  /* TG68K_FPU_Transcendental.vhd:572:73  */
  assign n11633 = n11561 ? x_cubed : n11627;
  /* TG68K_FPU_Transcendental.vhd:572:73  */
  assign n11634 = n11561 ? x_fifth : n11628;
  /* TG68K_FPU_Transcendental.vhd:572:73  */
  assign n11635 = n11561 ? x3_div6 : n11629;
  /* TG68K_FPU_Transcendental.vhd:572:73  */
  assign n11636 = n11561 ? x5_div120 : n11630;
  /* TG68K_FPU_Transcendental.vhd:602:108  */
  assign n11637 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:602:108  */
  assign n11639 = n11637 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:602:92  */
  assign n11640 = n11639[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:608:95  */
  assign n11641 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:608:111  */
  assign n11643 = $unsigned(n11641) > $unsigned(15'b100000000001001);
  /* TG68K_FPU_Transcendental.vhd:613:105  */
  assign n11644 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:614:106  */
  assign n11645 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:608:73  */
  assign n11647 = n11643 ? 15'b100000000001001 : n11644;
  /* TG68K_FPU_Transcendental.vhd:608:73  */
  assign n11649 = n11643 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n11645;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11651 = n11558 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11652 = n11558 ? result_sign : input_sign;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11653 = n11558 ? result_exp : n11647;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11654 = n11558 ? result_mant : n11649;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11655 = n11558 ? n11631 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11656 = n11558 ? n11640 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11658 = n11558 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11659 = n11561 & n11558;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11660 = n11558 ? n11633 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11661 = n11558 ? n11634 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11662 = n11558 ? n11635 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:570:65  */
  assign n11663 = n11558 ? n11636 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11664 = n11542 ? n11548 : n11651;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11665 = n11542 ? n11549 : n11652;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11666 = n11542 ? n11551 : n11653;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11667 = n11542 ? n11553 : n11654;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11668 = n11542 ? n11554 : n11655;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11669 = n11542 ? n11555 : n11656;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11670 = n11542 ? trans_inexact : n11658;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11671 = n11542 ? x_squared : n11632;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11672 = n11542 ? x_cubed : n11660;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11673 = n11542 ? x_fifth : n11661;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11674 = n11542 ? x3_div6 : n11662;
  /* TG68K_FPU_Transcendental.vhd:557:65  */
  assign n11675 = n11542 ? x5_div120 : n11663;
  /* TG68K_FPU_Transcendental.vhd:554:57  */
  assign n11677 = operation_code == 7'b0001111;
  /* TG68K_FPU_Transcendental.vhd:622:84  */
  assign n11678 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:622:84  */
  assign n11680 = n11678 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:632:116  */
  assign n11681 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:632:116  */
  assign n11683 = n11681 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:632:100  */
  assign n11684 = n11683[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:623:73  */
  assign n11686 = input_zero ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:623:73  */
  assign n11687 = input_zero ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:623:73  */
  assign n11689 = input_zero ? 15'b000000000000000 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:623:73  */
  assign n11691 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:623:73  */
  assign n11692 = input_zero ? series_sum : operand;
  /* TG68K_FPU_Transcendental.vhd:623:73  */
  assign n11693 = input_zero ? iteration_count : n11684;
  /* TG68K_FPU_Transcendental.vhd:634:87  */
  assign n11694 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:634:87  */
  assign n11696 = $signed(n11694) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU_Transcendental.vhd:636:92  */
  assign n11697 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:636:92  */
  assign n11699 = n11697 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:639:115  */
  assign n11700 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:639:152  */
  assign n11701 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:639:131  */
  assign n11702 = {32'b0, n11700};  //  uext
  /* TG68K_FPU_Transcendental.vhd:639:131  */
  assign n11703 = {32'b0, n11701};  //  uext
  /* TG68K_FPU_Transcendental.vhd:639:131  */
  assign n11704 = n11702 * n11703; // umul
  /* TG68K_FPU_Transcendental.vhd:639:89  */
  assign n11705 = {64'b0, n11704};  //  uext
  /* TG68K_FPU_Transcendental.vhd:641:95  */
  assign n11706 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:641:95  */
  assign n11708 = n11706 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:644:114  */
  assign n11709 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:644:152  */
  assign n11710 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:644:131  */
  assign n11711 = {32'b0, n11709};  //  uext
  /* TG68K_FPU_Transcendental.vhd:644:131  */
  assign n11712 = {32'b0, n11710};  //  uext
  /* TG68K_FPU_Transcendental.vhd:644:131  */
  assign n11713 = n11711 * n11712; // umul
  /* TG68K_FPU_Transcendental.vhd:644:89  */
  assign n11714 = {64'b0, n11713};  //  uext
  /* TG68K_FPU_Transcendental.vhd:646:95  */
  assign n11715 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:646:95  */
  assign n11717 = n11715 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:648:132  */
  assign n11718 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:648:149  */
  assign n11720 = n11718 / 32'b00000000000000000000000000000110; // udiv
  /* TG68K_FPU_Transcendental.vhd:648:109  */
  assign n11721 = {32'b0, n11720};  //  uext
  /* TG68K_FPU_Transcendental.vhd:649:95  */
  assign n11722 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:649:95  */
  assign n11724 = n11722 == 32'b00000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:652:89  */
  assign n11725 = {16'b0, x3_div6};  //  uext
  /* TG68K_FPU_Transcendental.vhd:651:133  */
  assign n11726 = series_sum + n11725;
  /* TG68K_FPU_Transcendental.vhd:653:95  */
  assign n11727 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:653:95  */
  assign n11729 = n11727 == 32'b00000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:656:112  */
  assign n11730 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:656:149  */
  assign n11731 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:656:129  */
  assign n11732 = {32'b0, n11730};  //  uext
  /* TG68K_FPU_Transcendental.vhd:656:129  */
  assign n11733 = {32'b0, n11731};  //  uext
  /* TG68K_FPU_Transcendental.vhd:656:129  */
  assign n11734 = n11732 * n11733; // umul
  /* TG68K_FPU_Transcendental.vhd:656:89  */
  assign n11735 = {64'b0, n11734};  //  uext
  /* TG68K_FPU_Transcendental.vhd:658:95  */
  assign n11736 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:658:95  */
  assign n11738 = n11736 == 32'b00000000000000000000000000000110;
  /* TG68K_FPU_Transcendental.vhd:660:139  */
  assign n11739 = x_fifth[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:660:111  */
  assign n11741 = n11739 >> 31'b0000000000000000000000000000111;
  /* TG68K_FPU_Transcendental.vhd:661:95  */
  assign n11742 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:661:95  */
  assign n11744 = n11742 == 32'b00000000000000000000000000000111;
  /* TG68K_FPU_Transcendental.vhd:664:89  */
  assign n11745 = {16'b0, x5_div120};  //  uext
  /* TG68K_FPU_Transcendental.vhd:663:133  */
  assign n11746 = series_sum + n11745;
  /* TG68K_FPU_Transcendental.vhd:661:73  */
  assign n11747 = n11744 ? n11746 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:658:73  */
  assign n11748 = n11738 ? series_sum : n11747;
  /* TG68K_FPU_Transcendental.vhd:658:73  */
  assign n11749 = n11738 ? n11741 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:653:73  */
  assign n11750 = n11729 ? series_sum : n11748;
  /* TG68K_FPU_Transcendental.vhd:653:73  */
  assign n11751 = n11729 ? n11735 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:653:73  */
  assign n11752 = n11729 ? x5_div120 : n11749;
  /* TG68K_FPU_Transcendental.vhd:649:73  */
  assign n11753 = n11724 ? n11726 : n11750;
  /* TG68K_FPU_Transcendental.vhd:649:73  */
  assign n11754 = n11724 ? x_fifth : n11751;
  /* TG68K_FPU_Transcendental.vhd:649:73  */
  assign n11755 = n11724 ? x5_div120 : n11752;
  /* TG68K_FPU_Transcendental.vhd:646:73  */
  assign n11756 = n11717 ? series_sum : n11753;
  /* TG68K_FPU_Transcendental.vhd:646:73  */
  assign n11757 = n11717 ? x_fifth : n11754;
  /* TG68K_FPU_Transcendental.vhd:646:73  */
  assign n11758 = n11717 ? n11721 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:646:73  */
  assign n11759 = n11717 ? x5_div120 : n11755;
  /* TG68K_FPU_Transcendental.vhd:641:73  */
  assign n11760 = n11708 ? series_sum : n11756;
  /* TG68K_FPU_Transcendental.vhd:641:73  */
  assign n11761 = n11708 ? n11714 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:641:73  */
  assign n11762 = n11708 ? x_fifth : n11757;
  /* TG68K_FPU_Transcendental.vhd:641:73  */
  assign n11763 = n11708 ? x3_div6 : n11758;
  /* TG68K_FPU_Transcendental.vhd:641:73  */
  assign n11764 = n11708 ? x5_div120 : n11759;
  /* TG68K_FPU_Transcendental.vhd:636:73  */
  assign n11765 = n11699 ? series_sum : n11760;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11766 = n11792 ? n11705 : x_squared;
  /* TG68K_FPU_Transcendental.vhd:636:73  */
  assign n11767 = n11699 ? x_cubed : n11761;
  /* TG68K_FPU_Transcendental.vhd:636:73  */
  assign n11768 = n11699 ? x_fifth : n11762;
  /* TG68K_FPU_Transcendental.vhd:636:73  */
  assign n11769 = n11699 ? x3_div6 : n11763;
  /* TG68K_FPU_Transcendental.vhd:636:73  */
  assign n11770 = n11699 ? x5_div120 : n11764;
  /* TG68K_FPU_Transcendental.vhd:666:108  */
  assign n11771 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:666:108  */
  assign n11773 = n11771 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:666:92  */
  assign n11774 = n11773[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:671:96  */
  assign n11776 = $unsigned(input_exp) >= $unsigned(15'b100000000000011);
  /* TG68K_FPU_Transcendental.vhd:673:132  */
  assign n11778 = input_exp + 15'b000000000000001;
  /* TG68K_FPU_Transcendental.vhd:677:105  */
  assign n11779 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:678:106  */
  assign n11780 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:671:73  */
  assign n11781 = n11776 ? n11778 : n11779;
  /* TG68K_FPU_Transcendental.vhd:671:73  */
  assign n11782 = n11776 ? input_mant : n11780;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11784 = n11696 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11785 = n11696 ? result_sign : input_sign;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11786 = n11696 ? result_exp : n11781;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11787 = n11696 ? result_mant : n11782;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11788 = n11696 ? n11765 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11789 = n11696 ? n11774 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11791 = n11696 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11792 = n11699 & n11696;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11793 = n11696 ? n11767 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11794 = n11696 ? n11768 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11795 = n11696 ? n11769 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:634:65  */
  assign n11796 = n11696 ? n11770 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11797 = n11680 ? n11686 : n11784;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11798 = n11680 ? n11687 : n11785;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11799 = n11680 ? n11689 : n11786;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11800 = n11680 ? n11691 : n11787;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11801 = n11680 ? n11692 : n11788;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11802 = n11680 ? n11693 : n11789;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11803 = n11680 ? trans_inexact : n11791;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11804 = n11680 ? x_squared : n11766;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11805 = n11680 ? x_cubed : n11793;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11806 = n11680 ? x_fifth : n11794;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11807 = n11680 ? x3_div6 : n11795;
  /* TG68K_FPU_Transcendental.vhd:622:65  */
  assign n11808 = n11680 ? x5_div120 : n11796;
  /* TG68K_FPU_Transcendental.vhd:619:57  */
  assign n11810 = operation_code == 7'b0001011;
  /* TG68K_FPU_Transcendental.vhd:686:84  */
  assign n11811 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:686:84  */
  assign n11813 = n11811 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:696:116  */
  assign n11814 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:696:116  */
  assign n11816 = n11814 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:696:100  */
  assign n11817 = n11816[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:687:73  */
  assign n11819 = input_zero ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:687:73  */
  assign n11821 = input_zero ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:687:73  */
  assign n11823 = input_zero ? 15'b011111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:687:73  */
  assign n11825 = input_zero ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:687:73  */
  assign n11827 = input_zero ? series_sum : 80'b00111111111111111000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:687:73  */
  assign n11828 = input_zero ? iteration_count : n11817;
  /* TG68K_FPU_Transcendental.vhd:698:87  */
  assign n11829 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:698:87  */
  assign n11831 = $signed(n11829) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU_Transcendental.vhd:700:92  */
  assign n11832 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:700:92  */
  assign n11834 = n11832 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:703:115  */
  assign n11835 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:703:152  */
  assign n11836 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:703:131  */
  assign n11837 = {32'b0, n11835};  //  uext
  /* TG68K_FPU_Transcendental.vhd:703:131  */
  assign n11838 = {32'b0, n11836};  //  uext
  /* TG68K_FPU_Transcendental.vhd:703:131  */
  assign n11839 = n11837 * n11838; // umul
  /* TG68K_FPU_Transcendental.vhd:703:89  */
  assign n11840 = {64'b0, n11839};  //  uext
  /* TG68K_FPU_Transcendental.vhd:705:95  */
  assign n11841 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:705:95  */
  assign n11843 = n11841 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:708:126  */
  assign n11844 = x_squared[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:708:96  */
  assign n11846 = n11844 >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:708:89  */
  assign n11847 = {16'b0, n11846};  //  uext
  /* TG68K_FPU_Transcendental.vhd:707:133  */
  assign n11848 = series_sum + n11847;
  /* TG68K_FPU_Transcendental.vhd:709:95  */
  assign n11849 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:709:95  */
  assign n11851 = n11849 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:712:114  */
  assign n11852 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:712:151  */
  assign n11853 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:712:131  */
  assign n11854 = {32'b0, n11852};  //  uext
  /* TG68K_FPU_Transcendental.vhd:712:131  */
  assign n11855 = {32'b0, n11853};  //  uext
  /* TG68K_FPU_Transcendental.vhd:712:131  */
  assign n11856 = n11854 * n11855; // umul
  /* TG68K_FPU_Transcendental.vhd:712:89  */
  assign n11857 = {64'b0, n11856};  //  uext
  /* TG68K_FPU_Transcendental.vhd:714:95  */
  assign n11858 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:714:95  */
  assign n11860 = n11858 == 32'b00000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:717:124  */
  assign n11861 = x_cubed[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:717:96  */
  assign n11863 = n11861 >> 31'b0000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:717:89  */
  assign n11864 = {16'b0, n11863};  //  uext
  /* TG68K_FPU_Transcendental.vhd:716:133  */
  assign n11865 = series_sum + n11864;
  /* TG68K_FPU_Transcendental.vhd:718:95  */
  assign n11866 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:718:95  */
  assign n11868 = n11866 == 32'b00000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:721:112  */
  assign n11869 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:721:149  */
  assign n11870 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:721:129  */
  assign n11871 = {32'b0, n11869};  //  uext
  /* TG68K_FPU_Transcendental.vhd:721:129  */
  assign n11872 = {32'b0, n11870};  //  uext
  /* TG68K_FPU_Transcendental.vhd:721:129  */
  assign n11873 = n11871 * n11872; // umul
  /* TG68K_FPU_Transcendental.vhd:721:89  */
  assign n11874 = {64'b0, n11873};  //  uext
  /* TG68K_FPU_Transcendental.vhd:723:95  */
  assign n11875 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:723:95  */
  assign n11877 = n11875 == 32'b00000000000000000000000000000110;
  /* TG68K_FPU_Transcendental.vhd:725:139  */
  assign n11878 = x_fifth[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:725:111  */
  assign n11880 = n11878 >> 31'b0000000000000000000000000001001;
  /* TG68K_FPU_Transcendental.vhd:726:95  */
  assign n11881 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:726:95  */
  assign n11883 = n11881 == 32'b00000000000000000000000000000111;
  /* TG68K_FPU_Transcendental.vhd:729:89  */
  assign n11884 = {16'b0, x5_div120};  //  uext
  /* TG68K_FPU_Transcendental.vhd:728:133  */
  assign n11885 = series_sum + n11884;
  /* TG68K_FPU_Transcendental.vhd:726:73  */
  assign n11886 = n11883 ? n11885 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:723:73  */
  assign n11887 = n11877 ? series_sum : n11886;
  /* TG68K_FPU_Transcendental.vhd:723:73  */
  assign n11888 = n11877 ? n11880 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:718:73  */
  assign n11889 = n11868 ? series_sum : n11887;
  /* TG68K_FPU_Transcendental.vhd:718:73  */
  assign n11890 = n11868 ? n11874 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:718:73  */
  assign n11891 = n11868 ? x5_div120 : n11888;
  /* TG68K_FPU_Transcendental.vhd:714:73  */
  assign n11892 = n11860 ? n11865 : n11889;
  /* TG68K_FPU_Transcendental.vhd:714:73  */
  assign n11893 = n11860 ? x_fifth : n11890;
  /* TG68K_FPU_Transcendental.vhd:714:73  */
  assign n11894 = n11860 ? x5_div120 : n11891;
  /* TG68K_FPU_Transcendental.vhd:709:73  */
  assign n11895 = n11851 ? series_sum : n11892;
  /* TG68K_FPU_Transcendental.vhd:709:73  */
  assign n11896 = n11851 ? n11857 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:709:73  */
  assign n11897 = n11851 ? x_fifth : n11893;
  /* TG68K_FPU_Transcendental.vhd:709:73  */
  assign n11898 = n11851 ? x5_div120 : n11894;
  /* TG68K_FPU_Transcendental.vhd:705:73  */
  assign n11899 = n11843 ? n11848 : n11895;
  /* TG68K_FPU_Transcendental.vhd:705:73  */
  assign n11900 = n11843 ? x_cubed : n11896;
  /* TG68K_FPU_Transcendental.vhd:705:73  */
  assign n11901 = n11843 ? x_fifth : n11897;
  /* TG68K_FPU_Transcendental.vhd:705:73  */
  assign n11902 = n11843 ? x5_div120 : n11898;
  /* TG68K_FPU_Transcendental.vhd:700:73  */
  assign n11903 = n11834 ? series_sum : n11899;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11904 = n11930 ? n11840 : x_squared;
  /* TG68K_FPU_Transcendental.vhd:700:73  */
  assign n11905 = n11834 ? x_cubed : n11900;
  /* TG68K_FPU_Transcendental.vhd:700:73  */
  assign n11906 = n11834 ? x_fifth : n11901;
  /* TG68K_FPU_Transcendental.vhd:700:73  */
  assign n11907 = n11834 ? x5_div120 : n11902;
  /* TG68K_FPU_Transcendental.vhd:731:108  */
  assign n11908 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:731:108  */
  assign n11910 = n11908 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:731:92  */
  assign n11911 = n11910[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:736:96  */
  assign n11913 = $unsigned(input_exp) >= $unsigned(15'b100000000000011);
  /* TG68K_FPU_Transcendental.vhd:738:132  */
  assign n11915 = input_exp + 15'b000000000000001;
  /* TG68K_FPU_Transcendental.vhd:742:105  */
  assign n11916 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:743:106  */
  assign n11917 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:736:73  */
  assign n11918 = n11913 ? n11915 : n11916;
  /* TG68K_FPU_Transcendental.vhd:736:73  */
  assign n11919 = n11913 ? input_mant : n11917;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11921 = n11831 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11923 = n11831 ? result_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11924 = n11831 ? result_exp : n11918;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11925 = n11831 ? result_mant : n11919;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11926 = n11831 ? n11903 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11927 = n11831 ? n11911 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11929 = n11831 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11930 = n11834 & n11831;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11931 = n11831 ? n11905 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11932 = n11831 ? n11906 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:698:65  */
  assign n11933 = n11831 ? n11907 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11934 = n11813 ? n11819 : n11921;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11935 = n11813 ? n11821 : n11923;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11936 = n11813 ? n11823 : n11924;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11937 = n11813 ? n11825 : n11925;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11938 = n11813 ? n11827 : n11926;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11939 = n11813 ? n11828 : n11927;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11940 = n11813 ? trans_inexact : n11929;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11941 = n11813 ? x_squared : n11904;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11942 = n11813 ? x_cubed : n11931;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11943 = n11813 ? x_fifth : n11932;
  /* TG68K_FPU_Transcendental.vhd:686:65  */
  assign n11944 = n11813 ? x5_div120 : n11933;
  /* TG68K_FPU_Transcendental.vhd:683:57  */
  assign n11946 = operation_code == 7'b0011001;
  /* TG68K_FPU_Transcendental.vhd:751:84  */
  assign n11947 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:751:84  */
  assign n11949 = n11947 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:760:104  */
  assign n11951 = $unsigned(input_exp) >= $unsigned(15'b100000000000010);
  /* TG68K_FPU_Transcendental.vhd:769:124  */
  assign n11952 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:769:124  */
  assign n11954 = n11952 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:769:108  */
  assign n11955 = n11954[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:760:81  */
  assign n11957 = n11951 ? 3'b110 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:760:81  */
  assign n11958 = n11951 ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:760:81  */
  assign n11960 = n11951 ? 15'b011111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:760:81  */
  assign n11962 = n11951 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:760:81  */
  assign n11963 = n11951 ? series_sum : operand;
  /* TG68K_FPU_Transcendental.vhd:760:81  */
  assign n11964 = n11951 ? iteration_count : n11955;
  /* TG68K_FPU_Transcendental.vhd:752:73  */
  assign n11966 = input_zero ? 3'b111 : n11957;
  /* TG68K_FPU_Transcendental.vhd:752:73  */
  assign n11967 = input_zero ? input_sign : n11958;
  /* TG68K_FPU_Transcendental.vhd:752:73  */
  assign n11969 = input_zero ? 15'b000000000000000 : n11960;
  /* TG68K_FPU_Transcendental.vhd:752:73  */
  assign n11971 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n11962;
  /* TG68K_FPU_Transcendental.vhd:752:73  */
  assign n11972 = input_zero ? series_sum : n11963;
  /* TG68K_FPU_Transcendental.vhd:752:73  */
  assign n11973 = input_zero ? iteration_count : n11964;
  /* TG68K_FPU_Transcendental.vhd:772:87  */
  assign n11974 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:772:87  */
  assign n11976 = $signed(n11974) <= $signed(32'b00000000000000000000000000001000);
  /* TG68K_FPU_Transcendental.vhd:775:92  */
  assign n11977 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:775:92  */
  assign n11979 = n11977 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:778:115  */
  assign n11980 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:778:152  */
  assign n11981 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:778:131  */
  assign n11982 = {32'b0, n11980};  //  uext
  /* TG68K_FPU_Transcendental.vhd:778:131  */
  assign n11983 = {32'b0, n11981};  //  uext
  /* TG68K_FPU_Transcendental.vhd:778:131  */
  assign n11984 = n11982 * n11983; // umul
  /* TG68K_FPU_Transcendental.vhd:778:89  */
  assign n11985 = {64'b0, n11984};  //  uext
  /* TG68K_FPU_Transcendental.vhd:780:95  */
  assign n11986 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:780:95  */
  assign n11988 = n11986 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:783:114  */
  assign n11989 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:783:152  */
  assign n11990 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:783:131  */
  assign n11991 = {32'b0, n11989};  //  uext
  /* TG68K_FPU_Transcendental.vhd:783:131  */
  assign n11992 = {32'b0, n11990};  //  uext
  /* TG68K_FPU_Transcendental.vhd:783:131  */
  assign n11993 = n11991 * n11992; // umul
  /* TG68K_FPU_Transcendental.vhd:783:89  */
  assign n11994 = {64'b0, n11993};  //  uext
  /* TG68K_FPU_Transcendental.vhd:785:95  */
  assign n11995 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:785:95  */
  assign n11997 = n11995 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:787:132  */
  assign n11998 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:787:149  */
  assign n12000 = n11998 / 32'b00000000000000000000000000000011; // udiv
  /* TG68K_FPU_Transcendental.vhd:787:109  */
  assign n12001 = {32'b0, n12000};  //  uext
  /* TG68K_FPU_Transcendental.vhd:788:95  */
  assign n12002 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:788:95  */
  assign n12004 = n12002 == 32'b00000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:791:89  */
  assign n12005 = {16'b0, x3_div6};  //  uext
  /* TG68K_FPU_Transcendental.vhd:790:133  */
  assign n12006 = series_sum - n12005;
  /* TG68K_FPU_Transcendental.vhd:792:95  */
  assign n12007 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:792:95  */
  assign n12009 = n12007 == 32'b00000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:795:112  */
  assign n12010 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:795:149  */
  assign n12011 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:795:129  */
  assign n12012 = {32'b0, n12010};  //  uext
  /* TG68K_FPU_Transcendental.vhd:795:129  */
  assign n12013 = {32'b0, n12011};  //  uext
  /* TG68K_FPU_Transcendental.vhd:795:129  */
  assign n12014 = n12012 * n12013; // umul
  /* TG68K_FPU_Transcendental.vhd:795:89  */
  assign n12015 = {64'b0, n12014};  //  uext
  /* TG68K_FPU_Transcendental.vhd:797:95  */
  assign n12016 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:797:95  */
  assign n12018 = n12016 == 32'b00000000000000000000000000000110;
  /* TG68K_FPU_Transcendental.vhd:799:146  */
  assign n12019 = x_fifth[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:799:163  */
  assign n12020 = {64'b0, n12019};  //  uext
  /* TG68K_FPU_Transcendental.vhd:799:163  */
  assign n12022 = $signed(n12020) * $signed(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010); // smul
  /* TG68K_FPU_Transcendental.vhd:799:118  */
  assign n12024 = n12022 >> 31'b0000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:799:111  */
  assign n12025 = n12024[63:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:800:95  */
  assign n12026 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:800:95  */
  assign n12028 = n12026 == 32'b00000000000000000000000000000111;
  /* TG68K_FPU_Transcendental.vhd:803:89  */
  assign n12029 = {16'b0, x5_div120};  //  uext
  /* TG68K_FPU_Transcendental.vhd:802:133  */
  assign n12030 = series_sum + n12029;
  /* TG68K_FPU_Transcendental.vhd:800:73  */
  assign n12031 = n12028 ? n12030 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:797:73  */
  assign n12032 = n12018 ? series_sum : n12031;
  /* TG68K_FPU_Transcendental.vhd:797:73  */
  assign n12033 = n12018 ? n12025 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:792:73  */
  assign n12034 = n12009 ? series_sum : n12032;
  /* TG68K_FPU_Transcendental.vhd:792:73  */
  assign n12035 = n12009 ? n12015 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:792:73  */
  assign n12036 = n12009 ? x5_div120 : n12033;
  /* TG68K_FPU_Transcendental.vhd:788:73  */
  assign n12037 = n12004 ? n12006 : n12034;
  /* TG68K_FPU_Transcendental.vhd:788:73  */
  assign n12038 = n12004 ? x_fifth : n12035;
  /* TG68K_FPU_Transcendental.vhd:788:73  */
  assign n12039 = n12004 ? x5_div120 : n12036;
  /* TG68K_FPU_Transcendental.vhd:785:73  */
  assign n12040 = n11997 ? series_sum : n12037;
  /* TG68K_FPU_Transcendental.vhd:785:73  */
  assign n12041 = n11997 ? x_fifth : n12038;
  /* TG68K_FPU_Transcendental.vhd:785:73  */
  assign n12042 = n11997 ? n12001 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:785:73  */
  assign n12043 = n11997 ? x5_div120 : n12039;
  /* TG68K_FPU_Transcendental.vhd:780:73  */
  assign n12044 = n11988 ? series_sum : n12040;
  /* TG68K_FPU_Transcendental.vhd:780:73  */
  assign n12045 = n11988 ? n11994 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:780:73  */
  assign n12046 = n11988 ? x_fifth : n12041;
  /* TG68K_FPU_Transcendental.vhd:780:73  */
  assign n12047 = n11988 ? x3_div6 : n12042;
  /* TG68K_FPU_Transcendental.vhd:780:73  */
  assign n12048 = n11988 ? x5_div120 : n12043;
  /* TG68K_FPU_Transcendental.vhd:775:73  */
  assign n12049 = n11979 ? series_sum : n12044;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12050 = n12077 ? n11985 : x_squared;
  /* TG68K_FPU_Transcendental.vhd:775:73  */
  assign n12051 = n11979 ? x_cubed : n12045;
  /* TG68K_FPU_Transcendental.vhd:775:73  */
  assign n12052 = n11979 ? x_fifth : n12046;
  /* TG68K_FPU_Transcendental.vhd:775:73  */
  assign n12053 = n11979 ? x3_div6 : n12047;
  /* TG68K_FPU_Transcendental.vhd:775:73  */
  assign n12054 = n11979 ? x5_div120 : n12048;
  /* TG68K_FPU_Transcendental.vhd:805:108  */
  assign n12055 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:805:108  */
  assign n12057 = n12055 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:805:92  */
  assign n12058 = n12057[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:811:95  */
  assign n12059 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:811:111  */
  assign n12061 = $unsigned(n12059) >= $unsigned(15'b011111111111111);
  /* TG68K_FPU_Transcendental.vhd:816:105  */
  assign n12062 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:817:106  */
  assign n12063 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:811:73  */
  assign n12065 = n12061 ? 15'b011111111111111 : n12062;
  /* TG68K_FPU_Transcendental.vhd:811:73  */
  assign n12067 = n12061 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n12063;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12069 = n11976 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12070 = n11976 ? result_sign : input_sign;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12071 = n11976 ? result_exp : n12065;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12072 = n11976 ? result_mant : n12067;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12073 = n11976 ? n12049 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12074 = n11976 ? n12058 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12076 = n11976 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12077 = n11979 & n11976;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12078 = n11976 ? n12051 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12079 = n11976 ? n12052 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12080 = n11976 ? n12053 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:772:65  */
  assign n12081 = n11976 ? n12054 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12082 = n11949 ? n11966 : n12069;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12083 = n11949 ? n11967 : n12070;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12084 = n11949 ? n11969 : n12071;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12085 = n11949 ? n11971 : n12072;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12086 = n11949 ? n11972 : n12073;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12087 = n11949 ? n11973 : n12074;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12088 = n11949 ? trans_inexact : n12076;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12089 = n11949 ? x_squared : n12050;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12090 = n11949 ? x_cubed : n12078;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12091 = n11949 ? x_fifth : n12079;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12092 = n11949 ? x3_div6 : n12080;
  /* TG68K_FPU_Transcendental.vhd:751:65  */
  assign n12093 = n11949 ? x5_div120 : n12081;
  /* TG68K_FPU_Transcendental.vhd:748:57  */
  assign n12095 = operation_code == 7'b0001001;
  /* TG68K_FPU_Transcendental.vhd:825:84  */
  assign n12096 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:825:84  */
  assign n12098 = n12096 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:827:96  */
  assign n12100 = $unsigned(input_exp) > $unsigned(15'b011111111111111);
  /* TG68K_FPU_Transcendental.vhd:828:97  */
  assign n12102 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:828:137  */
  assign n12104 = $unsigned(input_mant) > $unsigned(64'b1000000000000000000000000000000000000000000000000000000000000000);
  /* TG68K_FPU_Transcendental.vhd:828:122  */
  assign n12105 = n12104 & n12102;
  /* TG68K_FPU_Transcendental.vhd:827:121  */
  assign n12106 = n12100 | n12105;
  /* TG68K_FPU_Transcendental.vhd:841:99  */
  assign n12108 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:842:89  */
  assign n12109 = input_mant[63:62]; // extract
  /* TG68K_FPU_Transcendental.vhd:842:104  */
  assign n12111 = n12109 == 2'b10;
  /* TG68K_FPU_Transcendental.vhd:841:124  */
  assign n12112 = n12111 & n12108;
  /* TG68K_FPU_Transcendental.vhd:851:116  */
  assign n12113 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:851:116  */
  assign n12115 = n12113 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:851:100  */
  assign n12116 = n12115[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:841:73  */
  assign n12118 = n12112 ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:841:73  */
  assign n12119 = n12112 ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:841:73  */
  assign n12121 = n12112 ? 15'b011111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:841:73  */
  assign n12123 = n12112 ? 64'b1100100100001111110110101010001000100001011010001100001000110101 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:841:73  */
  assign n12124 = n12112 ? series_sum : operand;
  /* TG68K_FPU_Transcendental.vhd:841:73  */
  assign n12125 = n12112 ? iteration_count : n12116;
  /* TG68K_FPU_Transcendental.vhd:835:73  */
  assign n12127 = input_zero ? 3'b111 : n12118;
  /* TG68K_FPU_Transcendental.vhd:835:73  */
  assign n12128 = input_zero ? input_sign : n12119;
  /* TG68K_FPU_Transcendental.vhd:835:73  */
  assign n12130 = input_zero ? 15'b000000000000000 : n12121;
  /* TG68K_FPU_Transcendental.vhd:835:73  */
  assign n12132 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n12123;
  /* TG68K_FPU_Transcendental.vhd:835:73  */
  assign n12133 = input_zero ? series_sum : n12124;
  /* TG68K_FPU_Transcendental.vhd:835:73  */
  assign n12134 = input_zero ? iteration_count : n12125;
  /* TG68K_FPU_Transcendental.vhd:827:73  */
  assign n12136 = n12106 ? 3'b111 : n12127;
  /* TG68K_FPU_Transcendental.vhd:827:73  */
  assign n12138 = n12106 ? 1'b0 : n12128;
  /* TG68K_FPU_Transcendental.vhd:827:73  */
  assign n12140 = n12106 ? 15'b111111111111111 : n12130;
  /* TG68K_FPU_Transcendental.vhd:827:73  */
  assign n12142 = n12106 ? 64'b1100000000000000000000000000000000000000000000000000000000000000 : n12132;
  /* TG68K_FPU_Transcendental.vhd:827:73  */
  assign n12143 = n12106 ? series_sum : n12133;
  /* TG68K_FPU_Transcendental.vhd:827:73  */
  assign n12144 = n12106 ? iteration_count : n12134;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12146 = n12255 ? 1'b1 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:853:87  */
  assign n12147 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:853:87  */
  assign n12149 = $signed(n12147) <= $signed(32'b00000000000000000000000000001000);
  /* TG68K_FPU_Transcendental.vhd:855:92  */
  assign n12150 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:855:92  */
  assign n12152 = n12150 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:858:115  */
  assign n12153 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:858:152  */
  assign n12154 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:858:131  */
  assign n12155 = {32'b0, n12153};  //  uext
  /* TG68K_FPU_Transcendental.vhd:858:131  */
  assign n12156 = {32'b0, n12154};  //  uext
  /* TG68K_FPU_Transcendental.vhd:858:131  */
  assign n12157 = n12155 * n12156; // umul
  /* TG68K_FPU_Transcendental.vhd:858:89  */
  assign n12158 = {64'b0, n12157};  //  uext
  /* TG68K_FPU_Transcendental.vhd:860:95  */
  assign n12159 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:860:95  */
  assign n12161 = n12159 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:863:114  */
  assign n12162 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:863:152  */
  assign n12163 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:863:131  */
  assign n12164 = {32'b0, n12162};  //  uext
  /* TG68K_FPU_Transcendental.vhd:863:131  */
  assign n12165 = {32'b0, n12163};  //  uext
  /* TG68K_FPU_Transcendental.vhd:863:131  */
  assign n12166 = n12164 * n12165; // umul
  /* TG68K_FPU_Transcendental.vhd:863:89  */
  assign n12167 = {64'b0, n12166};  //  uext
  /* TG68K_FPU_Transcendental.vhd:865:95  */
  assign n12168 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:865:95  */
  assign n12170 = n12168 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:867:132  */
  assign n12171 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:867:149  */
  assign n12173 = n12171 / 32'b00000000000000000000000000000110; // udiv
  /* TG68K_FPU_Transcendental.vhd:867:109  */
  assign n12174 = {32'b0, n12173};  //  uext
  /* TG68K_FPU_Transcendental.vhd:868:95  */
  assign n12175 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:868:95  */
  assign n12177 = n12175 == 32'b00000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:871:89  */
  assign n12178 = {16'b0, x3_div6};  //  uext
  /* TG68K_FPU_Transcendental.vhd:870:133  */
  assign n12179 = series_sum + n12178;
  /* TG68K_FPU_Transcendental.vhd:872:95  */
  assign n12180 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:872:95  */
  assign n12182 = n12180 == 32'b00000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:875:112  */
  assign n12183 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:875:149  */
  assign n12184 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:875:129  */
  assign n12185 = {32'b0, n12183};  //  uext
  /* TG68K_FPU_Transcendental.vhd:875:129  */
  assign n12186 = {32'b0, n12184};  //  uext
  /* TG68K_FPU_Transcendental.vhd:875:129  */
  assign n12187 = n12185 * n12186; // umul
  /* TG68K_FPU_Transcendental.vhd:875:89  */
  assign n12188 = {64'b0, n12187};  //  uext
  /* TG68K_FPU_Transcendental.vhd:877:95  */
  assign n12189 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:877:95  */
  assign n12191 = n12189 == 32'b00000000000000000000000000000110;
  /* TG68K_FPU_Transcendental.vhd:879:146  */
  assign n12192 = x_fifth[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:879:163  */
  assign n12193 = {64'b0, n12192};  //  uext
  /* TG68K_FPU_Transcendental.vhd:879:163  */
  assign n12195 = $signed(n12193) * $signed(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011); // smul
  /* TG68K_FPU_Transcendental.vhd:879:118  */
  assign n12197 = n12195 >> 31'b0000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:879:111  */
  assign n12198 = n12197[63:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:880:95  */
  assign n12199 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:880:95  */
  assign n12201 = n12199 == 32'b00000000000000000000000000000111;
  /* TG68K_FPU_Transcendental.vhd:883:89  */
  assign n12202 = {16'b0, x5_div120};  //  uext
  /* TG68K_FPU_Transcendental.vhd:882:133  */
  assign n12203 = series_sum + n12202;
  /* TG68K_FPU_Transcendental.vhd:880:73  */
  assign n12204 = n12201 ? n12203 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:877:73  */
  assign n12205 = n12191 ? series_sum : n12204;
  /* TG68K_FPU_Transcendental.vhd:877:73  */
  assign n12206 = n12191 ? n12198 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:872:73  */
  assign n12207 = n12182 ? series_sum : n12205;
  /* TG68K_FPU_Transcendental.vhd:872:73  */
  assign n12208 = n12182 ? n12188 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:872:73  */
  assign n12209 = n12182 ? x5_div120 : n12206;
  /* TG68K_FPU_Transcendental.vhd:868:73  */
  assign n12210 = n12177 ? n12179 : n12207;
  /* TG68K_FPU_Transcendental.vhd:868:73  */
  assign n12211 = n12177 ? x_fifth : n12208;
  /* TG68K_FPU_Transcendental.vhd:868:73  */
  assign n12212 = n12177 ? x5_div120 : n12209;
  /* TG68K_FPU_Transcendental.vhd:865:73  */
  assign n12213 = n12170 ? series_sum : n12210;
  /* TG68K_FPU_Transcendental.vhd:865:73  */
  assign n12214 = n12170 ? x_fifth : n12211;
  /* TG68K_FPU_Transcendental.vhd:865:73  */
  assign n12215 = n12170 ? n12174 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:865:73  */
  assign n12216 = n12170 ? x5_div120 : n12212;
  /* TG68K_FPU_Transcendental.vhd:860:73  */
  assign n12217 = n12161 ? series_sum : n12213;
  /* TG68K_FPU_Transcendental.vhd:860:73  */
  assign n12218 = n12161 ? n12167 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:860:73  */
  assign n12219 = n12161 ? x_fifth : n12214;
  /* TG68K_FPU_Transcendental.vhd:860:73  */
  assign n12220 = n12161 ? x3_div6 : n12215;
  /* TG68K_FPU_Transcendental.vhd:860:73  */
  assign n12221 = n12161 ? x5_div120 : n12216;
  /* TG68K_FPU_Transcendental.vhd:855:73  */
  assign n12222 = n12152 ? series_sum : n12217;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12223 = n12243 ? n12158 : x_squared;
  /* TG68K_FPU_Transcendental.vhd:855:73  */
  assign n12224 = n12152 ? x_cubed : n12218;
  /* TG68K_FPU_Transcendental.vhd:855:73  */
  assign n12225 = n12152 ? x_fifth : n12219;
  /* TG68K_FPU_Transcendental.vhd:855:73  */
  assign n12226 = n12152 ? x3_div6 : n12220;
  /* TG68K_FPU_Transcendental.vhd:855:73  */
  assign n12227 = n12152 ? x5_div120 : n12221;
  /* TG68K_FPU_Transcendental.vhd:885:108  */
  assign n12228 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:885:108  */
  assign n12230 = n12228 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:885:92  */
  assign n12231 = n12230[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:890:97  */
  assign n12232 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:891:98  */
  assign n12233 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12235 = n12149 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12236 = n12149 ? result_sign : input_sign;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12237 = n12149 ? result_exp : n12232;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12238 = n12149 ? result_mant : n12233;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12239 = n12149 ? n12222 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12240 = n12149 ? n12231 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12242 = n12149 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12243 = n12152 & n12149;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12244 = n12149 ? n12224 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12245 = n12149 ? n12225 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12246 = n12149 ? n12226 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:853:65  */
  assign n12247 = n12149 ? n12227 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12248 = n12098 ? n12136 : n12235;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12249 = n12098 ? n12138 : n12236;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12250 = n12098 ? n12140 : n12237;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12251 = n12098 ? n12142 : n12238;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12252 = n12098 ? n12143 : n12239;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12253 = n12098 ? n12144 : n12240;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12254 = n12098 ? trans_inexact : n12242;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12255 = n12106 & n12098;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12256 = n12098 ? x_squared : n12223;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12257 = n12098 ? x_cubed : n12244;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12258 = n12098 ? x_fifth : n12245;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12259 = n12098 ? x3_div6 : n12246;
  /* TG68K_FPU_Transcendental.vhd:825:65  */
  assign n12260 = n12098 ? x5_div120 : n12247;
  /* TG68K_FPU_Transcendental.vhd:822:57  */
  assign n12262 = operation_code == 7'b0001100;
  /* TG68K_FPU_Transcendental.vhd:899:84  */
  assign n12263 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:899:84  */
  assign n12265 = n12263 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:901:96  */
  assign n12267 = $unsigned(input_exp) > $unsigned(15'b011111111111111);
  /* TG68K_FPU_Transcendental.vhd:902:97  */
  assign n12269 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:902:137  */
  assign n12271 = $unsigned(input_mant) > $unsigned(64'b1000000000000000000000000000000000000000000000000000000000000000);
  /* TG68K_FPU_Transcendental.vhd:902:122  */
  assign n12272 = n12271 & n12269;
  /* TG68K_FPU_Transcendental.vhd:901:121  */
  assign n12273 = n12267 | n12272;
  /* TG68K_FPU_Transcendental.vhd:915:99  */
  assign n12275 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:916:89  */
  assign n12276 = input_mant[63:62]; // extract
  /* TG68K_FPU_Transcendental.vhd:916:104  */
  assign n12278 = n12276 == 2'b10;
  /* TG68K_FPU_Transcendental.vhd:915:124  */
  assign n12279 = n12278 & n12275;
  /* TG68K_FPU_Transcendental.vhd:916:126  */
  assign n12280 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:916:111  */
  assign n12281 = n12280 & n12279;
  /* TG68K_FPU_Transcendental.vhd:922:99  */
  assign n12283 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:923:89  */
  assign n12284 = input_mant[63:62]; // extract
  /* TG68K_FPU_Transcendental.vhd:923:104  */
  assign n12286 = n12284 == 2'b10;
  /* TG68K_FPU_Transcendental.vhd:922:124  */
  assign n12287 = n12286 & n12283;
  /* TG68K_FPU_Transcendental.vhd:923:111  */
  assign n12288 = input_sign & n12287;
  /* TG68K_FPU_Transcendental.vhd:932:116  */
  assign n12289 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:932:116  */
  assign n12291 = n12289 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:932:100  */
  assign n12292 = n12291[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:922:73  */
  assign n12294 = n12288 ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:922:73  */
  assign n12296 = n12288 ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:922:73  */
  assign n12298 = n12288 ? 15'b100000000000000 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:922:73  */
  assign n12300 = n12288 ? 64'b1100100100001111110110101010001000100001011010001100001000110101 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:922:73  */
  assign n12302 = n12288 ? series_sum : 80'b00111111111111111100100100001111110110101010001000100001011010001100001000110101;
  /* TG68K_FPU_Transcendental.vhd:922:73  */
  assign n12303 = n12288 ? iteration_count : n12292;
  /* TG68K_FPU_Transcendental.vhd:915:73  */
  assign n12305 = n12281 ? 3'b111 : n12294;
  /* TG68K_FPU_Transcendental.vhd:915:73  */
  assign n12307 = n12281 ? 1'b0 : n12296;
  /* TG68K_FPU_Transcendental.vhd:915:73  */
  assign n12309 = n12281 ? 15'b000000000000000 : n12298;
  /* TG68K_FPU_Transcendental.vhd:915:73  */
  assign n12311 = n12281 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n12300;
  /* TG68K_FPU_Transcendental.vhd:915:73  */
  assign n12312 = n12281 ? series_sum : n12302;
  /* TG68K_FPU_Transcendental.vhd:915:73  */
  assign n12313 = n12281 ? iteration_count : n12303;
  /* TG68K_FPU_Transcendental.vhd:909:73  */
  assign n12315 = input_zero ? 3'b111 : n12305;
  /* TG68K_FPU_Transcendental.vhd:909:73  */
  assign n12317 = input_zero ? 1'b0 : n12307;
  /* TG68K_FPU_Transcendental.vhd:909:73  */
  assign n12319 = input_zero ? 15'b011111111111111 : n12309;
  /* TG68K_FPU_Transcendental.vhd:909:73  */
  assign n12321 = input_zero ? 64'b1100100100001111110110101010001000100001011010001100001000110101 : n12311;
  /* TG68K_FPU_Transcendental.vhd:909:73  */
  assign n12322 = input_zero ? series_sum : n12312;
  /* TG68K_FPU_Transcendental.vhd:909:73  */
  assign n12323 = input_zero ? iteration_count : n12313;
  /* TG68K_FPU_Transcendental.vhd:901:73  */
  assign n12325 = n12273 ? 3'b111 : n12315;
  /* TG68K_FPU_Transcendental.vhd:901:73  */
  assign n12327 = n12273 ? 1'b0 : n12317;
  /* TG68K_FPU_Transcendental.vhd:901:73  */
  assign n12329 = n12273 ? 15'b111111111111111 : n12319;
  /* TG68K_FPU_Transcendental.vhd:901:73  */
  assign n12331 = n12273 ? 64'b1100000000000000000000000000000000000000000000000000000000000000 : n12321;
  /* TG68K_FPU_Transcendental.vhd:901:73  */
  assign n12332 = n12273 ? series_sum : n12322;
  /* TG68K_FPU_Transcendental.vhd:901:73  */
  assign n12333 = n12273 ? iteration_count : n12323;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12335 = n12455 ? 1'b1 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:934:87  */
  assign n12336 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:934:87  */
  assign n12338 = $signed(n12336) <= $signed(32'b00000000000000000000000000001000);
  /* TG68K_FPU_Transcendental.vhd:937:92  */
  assign n12339 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:937:92  */
  assign n12341 = n12339 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:940:115  */
  assign n12342 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:940:152  */
  assign n12343 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:940:131  */
  assign n12344 = {32'b0, n12342};  //  uext
  /* TG68K_FPU_Transcendental.vhd:940:131  */
  assign n12345 = {32'b0, n12343};  //  uext
  /* TG68K_FPU_Transcendental.vhd:940:131  */
  assign n12346 = n12344 * n12345; // umul
  /* TG68K_FPU_Transcendental.vhd:940:89  */
  assign n12347 = {64'b0, n12346};  //  uext
  /* TG68K_FPU_Transcendental.vhd:942:95  */
  assign n12348 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:942:95  */
  assign n12350 = n12348 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:944:95  */
  assign n12351 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:945:138  */
  assign n12353 = 80'b00111111111111111100100100001111110110101010001000100001011010001100001000110101 - operand;
  /* TG68K_FPU_Transcendental.vhd:948:138  */
  assign n12355 = 80'b00111111111111111100100100001111110110101010001000100001011010001100001000110101 + operand;
  /* TG68K_FPU_Transcendental.vhd:944:81  */
  assign n12356 = n12351 ? n12353 : n12355;
  /* TG68K_FPU_Transcendental.vhd:951:95  */
  assign n12357 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:951:95  */
  assign n12359 = n12357 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:954:114  */
  assign n12360 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:954:152  */
  assign n12361 = input_mant[63:32]; // extract
  /* TG68K_FPU_Transcendental.vhd:954:131  */
  assign n12362 = {32'b0, n12360};  //  uext
  /* TG68K_FPU_Transcendental.vhd:954:131  */
  assign n12363 = {32'b0, n12361};  //  uext
  /* TG68K_FPU_Transcendental.vhd:954:131  */
  assign n12364 = n12362 * n12363; // umul
  /* TG68K_FPU_Transcendental.vhd:954:89  */
  assign n12365 = {64'b0, n12364};  //  uext
  /* TG68K_FPU_Transcendental.vhd:956:95  */
  assign n12366 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:956:95  */
  assign n12368 = n12366 == 32'b00000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:958:132  */
  assign n12369 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:958:149  */
  assign n12371 = n12369 / 32'b00000000000000000000000000000110; // udiv
  /* TG68K_FPU_Transcendental.vhd:958:109  */
  assign n12372 = {32'b0, n12371};  //  uext
  /* TG68K_FPU_Transcendental.vhd:959:95  */
  assign n12373 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:959:95  */
  assign n12375 = n12373 == 32'b00000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:961:95  */
  assign n12376 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:963:97  */
  assign n12377 = {16'b0, x3_div6};  //  uext
  /* TG68K_FPU_Transcendental.vhd:962:141  */
  assign n12378 = series_sum - n12377;
  /* TG68K_FPU_Transcendental.vhd:966:97  */
  assign n12379 = {16'b0, x3_div6};  //  uext
  /* TG68K_FPU_Transcendental.vhd:965:141  */
  assign n12380 = series_sum + n12379;
  /* TG68K_FPU_Transcendental.vhd:961:81  */
  assign n12381 = n12376 ? n12378 : n12380;
  /* TG68K_FPU_Transcendental.vhd:968:95  */
  assign n12382 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:968:95  */
  assign n12384 = n12382 == 32'b00000000000000000000000000000110;
  /* TG68K_FPU_Transcendental.vhd:971:112  */
  assign n12385 = x_cubed[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:971:149  */
  assign n12386 = x_squared[127:96]; // extract
  /* TG68K_FPU_Transcendental.vhd:971:129  */
  assign n12387 = {32'b0, n12385};  //  uext
  /* TG68K_FPU_Transcendental.vhd:971:129  */
  assign n12388 = {32'b0, n12386};  //  uext
  /* TG68K_FPU_Transcendental.vhd:971:129  */
  assign n12389 = n12387 * n12388; // umul
  /* TG68K_FPU_Transcendental.vhd:971:89  */
  assign n12390 = {64'b0, n12389};  //  uext
  /* TG68K_FPU_Transcendental.vhd:973:95  */
  assign n12391 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:973:95  */
  assign n12393 = n12391 == 32'b00000000000000000000000000000111;
  /* TG68K_FPU_Transcendental.vhd:975:146  */
  assign n12394 = x_fifth[127:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:975:163  */
  assign n12395 = {64'b0, n12394};  //  uext
  /* TG68K_FPU_Transcendental.vhd:975:163  */
  assign n12397 = $signed(n12395) * $signed(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011); // smul
  /* TG68K_FPU_Transcendental.vhd:975:118  */
  assign n12399 = n12397 >> 31'b0000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:975:111  */
  assign n12400 = n12399[63:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:973:73  */
  assign n12401 = n12393 ? n12400 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:968:73  */
  assign n12402 = n12384 ? n12390 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:968:73  */
  assign n12403 = n12384 ? x5_div120 : n12401;
  /* TG68K_FPU_Transcendental.vhd:959:73  */
  assign n12404 = n12375 ? n12381 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:959:73  */
  assign n12405 = n12375 ? x_fifth : n12402;
  /* TG68K_FPU_Transcendental.vhd:959:73  */
  assign n12406 = n12375 ? x5_div120 : n12403;
  /* TG68K_FPU_Transcendental.vhd:956:73  */
  assign n12407 = n12368 ? series_sum : n12404;
  /* TG68K_FPU_Transcendental.vhd:956:73  */
  assign n12408 = n12368 ? x_fifth : n12405;
  /* TG68K_FPU_Transcendental.vhd:956:73  */
  assign n12409 = n12368 ? n12372 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:956:73  */
  assign n12410 = n12368 ? x5_div120 : n12406;
  /* TG68K_FPU_Transcendental.vhd:951:73  */
  assign n12411 = n12359 ? series_sum : n12407;
  /* TG68K_FPU_Transcendental.vhd:951:73  */
  assign n12412 = n12359 ? n12365 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:951:73  */
  assign n12413 = n12359 ? x_fifth : n12408;
  /* TG68K_FPU_Transcendental.vhd:951:73  */
  assign n12414 = n12359 ? x3_div6 : n12409;
  /* TG68K_FPU_Transcendental.vhd:951:73  */
  assign n12415 = n12359 ? x5_div120 : n12410;
  /* TG68K_FPU_Transcendental.vhd:942:73  */
  assign n12416 = n12350 ? n12356 : n12411;
  /* TG68K_FPU_Transcendental.vhd:942:73  */
  assign n12417 = n12350 ? x_cubed : n12412;
  /* TG68K_FPU_Transcendental.vhd:942:73  */
  assign n12418 = n12350 ? x_fifth : n12413;
  /* TG68K_FPU_Transcendental.vhd:942:73  */
  assign n12419 = n12350 ? x3_div6 : n12414;
  /* TG68K_FPU_Transcendental.vhd:942:73  */
  assign n12420 = n12350 ? x5_div120 : n12415;
  /* TG68K_FPU_Transcendental.vhd:937:73  */
  assign n12421 = n12341 ? series_sum : n12416;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12422 = n12443 ? n12347 : x_squared;
  /* TG68K_FPU_Transcendental.vhd:937:73  */
  assign n12423 = n12341 ? x_cubed : n12417;
  /* TG68K_FPU_Transcendental.vhd:937:73  */
  assign n12424 = n12341 ? x_fifth : n12418;
  /* TG68K_FPU_Transcendental.vhd:937:73  */
  assign n12425 = n12341 ? x3_div6 : n12419;
  /* TG68K_FPU_Transcendental.vhd:937:73  */
  assign n12426 = n12341 ? x5_div120 : n12420;
  /* TG68K_FPU_Transcendental.vhd:977:108  */
  assign n12427 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:977:108  */
  assign n12429 = n12427 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:977:92  */
  assign n12430 = n12429[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:982:97  */
  assign n12431 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:983:98  */
  assign n12432 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12434 = n12338 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12436 = n12338 ? result_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12437 = n12338 ? result_exp : n12431;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12438 = n12338 ? result_mant : n12432;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12439 = n12338 ? n12421 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12440 = n12338 ? n12430 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12442 = n12338 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12443 = n12341 & n12338;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12444 = n12338 ? n12423 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12445 = n12338 ? n12424 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12446 = n12338 ? n12425 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:934:65  */
  assign n12447 = n12338 ? n12426 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12448 = n12265 ? n12325 : n12434;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12449 = n12265 ? n12327 : n12436;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12450 = n12265 ? n12329 : n12437;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12451 = n12265 ? n12331 : n12438;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12452 = n12265 ? n12332 : n12439;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12453 = n12265 ? n12333 : n12440;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12454 = n12265 ? trans_inexact : n12442;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12455 = n12273 & n12265;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12456 = n12265 ? x_squared : n12422;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12457 = n12265 ? x_cubed : n12444;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12458 = n12265 ? x_fifth : n12445;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12459 = n12265 ? x3_div6 : n12446;
  /* TG68K_FPU_Transcendental.vhd:899:65  */
  assign n12460 = n12265 ? x5_div120 : n12447;
  /* TG68K_FPU_Transcendental.vhd:895:57  */
  assign n12462 = operation_code == 7'b0011100;
  /* TG68K_FPU_Transcendental.vhd:995:91  */
  assign n12464 = $unsigned(input_exp) < $unsigned(15'b011111111110101);
  /* TG68K_FPU_Transcendental.vhd:995:65  */
  assign n12467 = n12464 ? 3'b110 : 3'b101;
  /* TG68K_FPU_Transcendental.vhd:995:65  */
  assign n12469 = n12464 ? cordic_iteration : 5'b00000;
  /* TG68K_FPU_Transcendental.vhd:995:65  */
  assign n12470 = n12464 ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:995:65  */
  assign n12471 = n12464 ? input_exp : result_exp;
  /* TG68K_FPU_Transcendental.vhd:995:65  */
  assign n12472 = n12464 ? input_mant : result_mant;
  /* TG68K_FPU_Transcendental.vhd:989:65  */
  assign n12474 = input_zero ? 3'b111 : n12467;
  /* TG68K_FPU_Transcendental.vhd:989:65  */
  assign n12475 = input_zero ? cordic_iteration : n12469;
  /* TG68K_FPU_Transcendental.vhd:989:65  */
  assign n12476 = input_zero ? input_sign : n12470;
  /* TG68K_FPU_Transcendental.vhd:989:65  */
  assign n12478 = input_zero ? 15'b000000000000000 : n12471;
  /* TG68K_FPU_Transcendental.vhd:989:65  */
  assign n12480 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n12472;
  /* TG68K_FPU_Transcendental.vhd:987:57  */
  assign n12482 = operation_code == 7'b0001010;
  /* TG68K_FPU_Transcendental.vhd:1009:84  */
  assign n12483 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1009:84  */
  assign n12485 = n12483 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1011:96  */
  assign n12487 = $unsigned(input_exp) >= $unsigned(15'b011111111111111);
  /* TG68K_FPU_Transcendental.vhd:1025:116  */
  assign n12488 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1025:116  */
  assign n12490 = n12488 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1025:100  */
  assign n12491 = n12490[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1018:73  */
  assign n12493 = input_zero ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:1018:73  */
  assign n12494 = input_zero ? input_sign : result_sign;
  /* TG68K_FPU_Transcendental.vhd:1018:73  */
  assign n12496 = input_zero ? 15'b000000000000000 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:1018:73  */
  assign n12498 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:1018:73  */
  assign n12499 = input_zero ? iteration_count : n12491;
  /* TG68K_FPU_Transcendental.vhd:1011:73  */
  assign n12501 = n12487 ? 3'b111 : n12493;
  /* TG68K_FPU_Transcendental.vhd:1011:73  */
  assign n12503 = n12487 ? 1'b0 : n12494;
  /* TG68K_FPU_Transcendental.vhd:1011:73  */
  assign n12505 = n12487 ? 15'b111111111111111 : n12496;
  /* TG68K_FPU_Transcendental.vhd:1011:73  */
  assign n12507 = n12487 ? 64'b1100000000000000000000000000000000000000000000000000000000000000 : n12498;
  /* TG68K_FPU_Transcendental.vhd:1011:73  */
  assign n12508 = n12487 ? iteration_count : n12499;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12510 = n12531 ? 1'b1 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:1027:87  */
  assign n12511 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1027:87  */
  assign n12513 = $signed(n12511) < $signed(32'b00000000000000000000000000000110);
  /* TG68K_FPU_Transcendental.vhd:1028:108  */
  assign n12514 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1028:108  */
  assign n12516 = n12514 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1028:92  */
  assign n12517 = n12516[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1027:65  */
  assign n12519 = n12513 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1027:65  */
  assign n12520 = n12513 ? result_sign : input_sign;
  /* TG68K_FPU_Transcendental.vhd:1027:65  */
  assign n12521 = n12513 ? result_exp : input_exp;
  /* TG68K_FPU_Transcendental.vhd:1027:65  */
  assign n12522 = n12513 ? result_mant : input_mant;
  /* TG68K_FPU_Transcendental.vhd:1027:65  */
  assign n12523 = n12513 ? n12517 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12524 = n12485 ? n12501 : n12519;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12525 = n12485 ? n12503 : n12520;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12526 = n12485 ? n12505 : n12521;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12527 = n12485 ? n12507 : n12522;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12528 = n12485 ? n12508 : n12523;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12530 = n12485 ? trans_inexact : 1'b1;
  /* TG68K_FPU_Transcendental.vhd:1009:65  */
  assign n12531 = n12487 & n12485;
  /* TG68K_FPU_Transcendental.vhd:1007:57  */
  assign n12533 = operation_code == 7'b0001101;
  /* TG68K_FPU_Transcendental.vhd:1042:84  */
  assign n12534 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1042:84  */
  assign n12536 = n12534 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1051:125  */
  assign n12538 = $unsigned(input_exp) > $unsigned(15'b100000000000101);
  /* TG68K_FPU_Transcendental.vhd:1051:101  */
  assign n12539 = n12538 & input_sign;
  /* TG68K_FPU_Transcendental.vhd:1058:98  */
  assign n12540 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:1058:128  */
  assign n12542 = $unsigned(input_exp) > $unsigned(15'b100000000000101);
  /* TG68K_FPU_Transcendental.vhd:1058:104  */
  assign n12543 = n12542 & n12540;
  /* TG68K_FPU_Transcendental.vhd:1070:124  */
  assign n12544 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1070:124  */
  assign n12546 = n12544 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1070:108  */
  assign n12547 = n12546[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12549 = n12543 ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12551 = n12543 ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12553 = n12543 ? 15'b111111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12555 = n12543 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12557 = n12543 ? series_term : 80'b00111111111111111000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12559 = n12543 ? series_sum : 80'b00111111111111111000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12560 = n12543 ? iteration_count : n12547;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12562 = n12543 ? 1'b1 : trans_overflow;
  /* TG68K_FPU_Transcendental.vhd:1058:81  */
  assign n12563 = n12543 ? exp_argument : operand;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12565 = n12539 ? 3'b111 : n12549;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12567 = n12539 ? 1'b0 : n12551;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12569 = n12539 ? 15'b000000000000000 : n12553;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12571 = n12539 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n12555;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12572 = n12539 ? series_term : n12557;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12573 = n12539 ? series_sum : n12559;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12574 = n12539 ? iteration_count : n12560;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12575 = n12539 ? trans_overflow : n12562;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12577 = n12539 ? 1'b1 : trans_underflow;
  /* TG68K_FPU_Transcendental.vhd:1051:81  */
  assign n12578 = n12539 ? exp_argument : n12563;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12580 = input_zero ? 3'b111 : n12565;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12582 = input_zero ? 1'b0 : n12567;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12584 = input_zero ? 15'b011111111111111 : n12569;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12586 = input_zero ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n12571;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12587 = input_zero ? series_term : n12572;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12588 = input_zero ? series_sum : n12573;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12589 = input_zero ? iteration_count : n12574;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12590 = input_zero ? trans_overflow : n12575;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12591 = input_zero ? trans_underflow : n12577;
  /* TG68K_FPU_Transcendental.vhd:1043:73  */
  assign n12592 = input_zero ? exp_argument : n12578;
  /* TG68K_FPU_Transcendental.vhd:1073:87  */
  assign n12593 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1073:87  */
  assign n12595 = $signed(n12593) <= $signed(32'b00000000000000000000000000000110);
  /* TG68K_FPU_Transcendental.vhd:1075:92  */
  assign n12596 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1075:92  */
  assign n12598 = n12596 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1078:133  */
  assign n12599 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1079:95  */
  assign n12600 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1079:95  */
  assign n12602 = n12600 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:1082:117  */
  assign n12603 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1082:156  */
  assign n12604 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1082:133  */
  assign n12605 = {16'b0, n12603};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1082:133  */
  assign n12606 = {16'b0, n12604};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1082:133  */
  assign n12607 = n12605 * n12606; // umul
  /* TG68K_FPU_Transcendental.vhd:1082:172  */
  assign n12609 = n12607 / 32'b00000000000000000000000000000010; // udiv
  /* TG68K_FPU_Transcendental.vhd:1082:89  */
  assign n12610 = {48'b0, n12609};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1084:133  */
  assign n12611 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1085:95  */
  assign n12612 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1085:95  */
  assign n12614 = n12612 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:1088:117  */
  assign n12615 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1088:156  */
  assign n12616 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1088:133  */
  assign n12617 = {16'b0, n12615};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1088:133  */
  assign n12618 = {16'b0, n12616};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1088:133  */
  assign n12619 = n12617 * n12618; // umul
  /* TG68K_FPU_Transcendental.vhd:1089:117  */
  assign n12620 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1088:172  */
  assign n12621 = {16'b0, n12619};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1088:172  */
  assign n12622 = {32'b0, n12620};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1088:172  */
  assign n12623 = n12621 * n12622; // umul
  /* TG68K_FPU_Transcendental.vhd:1089:133  */
  assign n12625 = n12623 / 48'b000000000000000000000000000000000000000000000110; // udiv
  /* TG68K_FPU_Transcendental.vhd:1088:89  */
  assign n12626 = {32'b0, n12625};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1091:133  */
  assign n12627 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1092:95  */
  assign n12628 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1092:95  */
  assign n12630 = n12628 == 32'b00000000000000000000000000000100;
  /* TG68K_FPU_Transcendental.vhd:1095:89  */
  assign n12632 = exp_argument >> 31'b0000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:1097:133  */
  assign n12633 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1092:73  */
  assign n12634 = n12630 ? n12632 : series_term;
  /* TG68K_FPU_Transcendental.vhd:1092:73  */
  assign n12635 = n12630 ? n12633 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:1085:73  */
  assign n12636 = n12614 ? n12626 : n12634;
  /* TG68K_FPU_Transcendental.vhd:1085:73  */
  assign n12637 = n12614 ? n12627 : n12635;
  /* TG68K_FPU_Transcendental.vhd:1079:73  */
  assign n12638 = n12602 ? n12610 : n12636;
  /* TG68K_FPU_Transcendental.vhd:1079:73  */
  assign n12639 = n12602 ? n12611 : n12637;
  /* TG68K_FPU_Transcendental.vhd:1075:73  */
  assign n12640 = n12598 ? exp_argument : n12638;
  /* TG68K_FPU_Transcendental.vhd:1075:73  */
  assign n12641 = n12598 ? n12599 : n12639;
  /* TG68K_FPU_Transcendental.vhd:1102:108  */
  assign n12642 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1102:108  */
  assign n12644 = n12642 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1102:92  */
  assign n12645 = n12644[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1106:98  */
  assign n12646 = series_sum[79]; // extract
  /* TG68K_FPU_Transcendental.vhd:1107:97  */
  assign n12647 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:1108:98  */
  assign n12648 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12650 = n12595 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12651 = n12595 ? result_sign : n12646;
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12652 = n12595 ? result_exp : n12647;
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12653 = n12595 ? result_mant : n12648;
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12654 = n12595 ? n12640 : series_term;
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12655 = n12595 ? n12641 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12656 = n12595 ? n12645 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:1073:65  */
  assign n12658 = n12595 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12659 = n12536 ? n12580 : n12650;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12660 = n12536 ? n12582 : n12651;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12661 = n12536 ? n12584 : n12652;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12662 = n12536 ? n12586 : n12653;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12663 = n12536 ? n12587 : n12654;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12664 = n12536 ? n12588 : n12655;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12665 = n12536 ? n12589 : n12656;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12666 = n12536 ? n12590 : trans_overflow;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12667 = n12536 ? n12591 : trans_underflow;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12668 = n12536 ? trans_inexact : n12658;
  /* TG68K_FPU_Transcendental.vhd:1042:65  */
  assign n12669 = n12536 ? n12592 : exp_argument;
  /* TG68K_FPU_Transcendental.vhd:1040:57  */
  assign n12671 = operation_code == 7'b0010000;
  /* TG68K_FPU_Transcendental.vhd:1114:84  */
  assign n12672 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1114:84  */
  assign n12674 = n12672 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1123:125  */
  assign n12676 = $unsigned(input_exp) > $unsigned(15'b100000000000101);
  /* TG68K_FPU_Transcendental.vhd:1123:101  */
  assign n12677 = n12676 & input_sign;
  /* TG68K_FPU_Transcendental.vhd:1130:98  */
  assign n12678 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:1130:128  */
  assign n12680 = $unsigned(input_exp) > $unsigned(15'b100000000000101);
  /* TG68K_FPU_Transcendental.vhd:1130:104  */
  assign n12681 = n12680 & n12678;
  /* TG68K_FPU_Transcendental.vhd:1142:124  */
  assign n12682 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1142:124  */
  assign n12684 = n12682 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1142:108  */
  assign n12685 = n12684[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12687 = n12681 ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12689 = n12681 ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12691 = n12681 ? 15'b111111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12693 = n12681 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12694 = n12681 ? series_term : operand;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12695 = n12681 ? series_sum : operand;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12696 = n12681 ? iteration_count : n12685;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12698 = n12681 ? 1'b1 : trans_overflow;
  /* TG68K_FPU_Transcendental.vhd:1130:81  */
  assign n12699 = n12681 ? exp_argument : operand;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12701 = n12677 ? 3'b111 : n12687;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12703 = n12677 ? 1'b1 : n12689;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12705 = n12677 ? 15'b011111111111111 : n12691;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12707 = n12677 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n12693;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12708 = n12677 ? series_term : n12694;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12709 = n12677 ? series_sum : n12695;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12710 = n12677 ? iteration_count : n12696;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12711 = n12677 ? trans_overflow : n12698;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12713 = n12677 ? 1'b1 : trans_underflow;
  /* TG68K_FPU_Transcendental.vhd:1123:81  */
  assign n12714 = n12677 ? exp_argument : n12699;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12716 = input_zero ? 3'b111 : n12701;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12718 = input_zero ? 1'b0 : n12703;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12720 = input_zero ? 15'b000000000000000 : n12705;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12722 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n12707;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12723 = input_zero ? series_term : n12708;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12724 = input_zero ? series_sum : n12709;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12725 = input_zero ? iteration_count : n12710;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12726 = input_zero ? trans_overflow : n12711;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12727 = input_zero ? trans_underflow : n12713;
  /* TG68K_FPU_Transcendental.vhd:1115:73  */
  assign n12728 = input_zero ? exp_argument : n12714;
  /* TG68K_FPU_Transcendental.vhd:1145:87  */
  assign n12729 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1145:87  */
  assign n12731 = $signed(n12729) <= $signed(32'b00000000000000000000000000000101);
  /* TG68K_FPU_Transcendental.vhd:1147:92  */
  assign n12732 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1147:92  */
  assign n12734 = n12732 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1150:117  */
  assign n12735 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1150:156  */
  assign n12736 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1150:133  */
  assign n12737 = {16'b0, n12735};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1150:133  */
  assign n12738 = {16'b0, n12736};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1150:133  */
  assign n12739 = n12737 * n12738; // umul
  /* TG68K_FPU_Transcendental.vhd:1150:172  */
  assign n12741 = n12739 / 32'b00000000000000000000000000000010; // udiv
  /* TG68K_FPU_Transcendental.vhd:1150:89  */
  assign n12742 = {48'b0, n12741};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1152:133  */
  assign n12743 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1153:95  */
  assign n12744 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1153:95  */
  assign n12746 = n12744 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:1156:117  */
  assign n12747 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1156:156  */
  assign n12748 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1156:133  */
  assign n12749 = {16'b0, n12747};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1156:133  */
  assign n12750 = {16'b0, n12748};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1156:133  */
  assign n12751 = n12749 * n12750; // umul
  /* TG68K_FPU_Transcendental.vhd:1157:117  */
  assign n12752 = exp_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1156:172  */
  assign n12753 = {16'b0, n12751};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1156:172  */
  assign n12754 = {32'b0, n12752};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1156:172  */
  assign n12755 = n12753 * n12754; // umul
  /* TG68K_FPU_Transcendental.vhd:1157:133  */
  assign n12757 = n12755 / 48'b000000000000000000000000000000000000000000000110; // udiv
  /* TG68K_FPU_Transcendental.vhd:1156:89  */
  assign n12758 = {32'b0, n12757};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1159:133  */
  assign n12759 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1160:95  */
  assign n12760 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1160:95  */
  assign n12762 = n12760 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:1163:89  */
  assign n12764 = exp_argument >> 31'b0000000000000000000000000000101;
  /* TG68K_FPU_Transcendental.vhd:1165:133  */
  assign n12765 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1160:73  */
  assign n12766 = n12762 ? n12764 : series_term;
  /* TG68K_FPU_Transcendental.vhd:1160:73  */
  assign n12767 = n12762 ? n12765 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:1153:73  */
  assign n12768 = n12746 ? n12758 : n12766;
  /* TG68K_FPU_Transcendental.vhd:1153:73  */
  assign n12769 = n12746 ? n12759 : n12767;
  /* TG68K_FPU_Transcendental.vhd:1147:73  */
  assign n12770 = n12734 ? n12742 : n12768;
  /* TG68K_FPU_Transcendental.vhd:1147:73  */
  assign n12771 = n12734 ? n12743 : n12769;
  /* TG68K_FPU_Transcendental.vhd:1170:108  */
  assign n12772 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1170:108  */
  assign n12774 = n12772 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1170:92  */
  assign n12775 = n12774[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1174:98  */
  assign n12776 = series_sum[79]; // extract
  /* TG68K_FPU_Transcendental.vhd:1175:97  */
  assign n12777 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:1176:98  */
  assign n12778 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12780 = n12731 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12781 = n12731 ? result_sign : n12776;
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12782 = n12731 ? result_exp : n12777;
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12783 = n12731 ? result_mant : n12778;
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12784 = n12731 ? n12770 : series_term;
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12785 = n12731 ? n12771 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12786 = n12731 ? n12775 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:1145:65  */
  assign n12788 = n12731 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12789 = n12674 ? n12716 : n12780;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12790 = n12674 ? n12718 : n12781;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12791 = n12674 ? n12720 : n12782;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12792 = n12674 ? n12722 : n12783;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12793 = n12674 ? n12723 : n12784;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12794 = n12674 ? n12724 : n12785;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12795 = n12674 ? n12725 : n12786;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12796 = n12674 ? n12726 : trans_overflow;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12797 = n12674 ? n12727 : trans_underflow;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12798 = n12674 ? trans_inexact : n12788;
  /* TG68K_FPU_Transcendental.vhd:1114:65  */
  assign n12799 = n12674 ? n12728 : exp_argument;
  /* TG68K_FPU_Transcendental.vhd:1112:57  */
  assign n12801 = operation_code == 7'b0000111;
  /* TG68K_FPU_Transcendental.vhd:1182:84  */
  assign n12802 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1182:84  */
  assign n12804 = n12802 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1183:117  */
  assign n12806 = $unsigned(input_exp) >= $unsigned(15'b011111111111111);
  /* TG68K_FPU_Transcendental.vhd:1183:93  */
  assign n12807 = n12806 & input_sign;
  /* TG68K_FPU_Transcendental.vhd:1196:99  */
  assign n12809 = input_exp == 15'b011111111111111;
  /* TG68K_FPU_Transcendental.vhd:1197:90  */
  assign n12811 = input_mant == 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1196:124  */
  assign n12812 = n12811 & n12809;
  /* TG68K_FPU_Transcendental.vhd:1197:112  */
  assign n12813 = input_sign & n12812;
  /* TG68K_FPU_Transcendental.vhd:1209:116  */
  assign n12814 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1209:116  */
  assign n12816 = n12814 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1209:100  */
  assign n12817 = n12816[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12819 = n12813 ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12821 = n12813 ? 1'b1 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12823 = n12813 ? 15'b111111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12825 = n12813 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12826 = n12813 ? series_term : operand;
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12827 = n12813 ? series_sum : operand;
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12828 = n12813 ? iteration_count : n12817;
  /* TG68K_FPU_Transcendental.vhd:1196:73  */
  assign n12829 = n12813 ? log_argument : operand;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12831 = input_zero ? 3'b111 : n12819;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12833 = input_zero ? 1'b0 : n12821;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12835 = input_zero ? 15'b000000000000000 : n12823;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12837 = input_zero ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n12825;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12838 = input_zero ? series_term : n12826;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12839 = input_zero ? series_sum : n12827;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12840 = input_zero ? iteration_count : n12828;
  /* TG68K_FPU_Transcendental.vhd:1190:73  */
  assign n12841 = input_zero ? log_argument : n12829;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12843 = n12807 ? 3'b111 : n12831;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12845 = n12807 ? 1'b0 : n12833;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12847 = n12807 ? 15'b111111111111111 : n12835;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12849 = n12807 ? 64'b1100000000000000000000000000000000000000000000000000000000000000 : n12837;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12850 = n12807 ? series_term : n12838;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12851 = n12807 ? series_sum : n12839;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12852 = n12807 ? iteration_count : n12840;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12854 = n12930 ? 1'b1 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:1183:73  */
  assign n12855 = n12807 ? log_argument : n12841;
  /* TG68K_FPU_Transcendental.vhd:1211:87  */
  assign n12856 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1211:87  */
  assign n12858 = $signed(n12856) <= $signed(32'b00000000000000000000000000000101);
  /* TG68K_FPU_Transcendental.vhd:1213:92  */
  assign n12859 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1213:92  */
  assign n12861 = n12859 == 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1216:117  */
  assign n12862 = log_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1216:156  */
  assign n12863 = log_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1216:133  */
  assign n12864 = {16'b0, n12862};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1216:133  */
  assign n12865 = {16'b0, n12863};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1216:133  */
  assign n12866 = n12864 * n12865; // umul
  /* TG68K_FPU_Transcendental.vhd:1216:172  */
  assign n12868 = n12866 / 32'b00000000000000000000000000000010; // udiv
  /* TG68K_FPU_Transcendental.vhd:1216:89  */
  assign n12869 = {48'b0, n12868};  //  uext
  assign n12871 = n12869[78:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1219:133  */
  assign n12872 = series_sum - series_term;
  /* TG68K_FPU_Transcendental.vhd:1220:95  */
  assign n12873 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1220:95  */
  assign n12875 = n12873 == 32'b00000000000000000000000000000010;
  /* TG68K_FPU_Transcendental.vhd:1223:117  */
  assign n12876 = log_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1223:156  */
  assign n12877 = log_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1223:133  */
  assign n12878 = {16'b0, n12876};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1223:133  */
  assign n12879 = {16'b0, n12877};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1223:133  */
  assign n12880 = n12878 * n12879; // umul
  /* TG68K_FPU_Transcendental.vhd:1224:117  */
  assign n12881 = log_argument[63:48]; // extract
  /* TG68K_FPU_Transcendental.vhd:1223:172  */
  assign n12882 = {16'b0, n12880};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1223:172  */
  assign n12883 = {32'b0, n12881};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1223:172  */
  assign n12884 = n12882 * n12883; // umul
  /* TG68K_FPU_Transcendental.vhd:1224:133  */
  assign n12886 = n12884 / 48'b000000000000000000000000000000000000000000000011; // udiv
  /* TG68K_FPU_Transcendental.vhd:1223:89  */
  assign n12887 = {32'b0, n12886};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1226:133  */
  assign n12888 = series_sum + series_term;
  /* TG68K_FPU_Transcendental.vhd:1227:95  */
  assign n12889 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1227:95  */
  assign n12891 = n12889 == 32'b00000000000000000000000000000011;
  /* TG68K_FPU_Transcendental.vhd:1230:89  */
  assign n12893 = log_argument >> 31'b0000000000000000000000000000010;
  assign n12895 = n12893[78:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1233:133  */
  assign n12896 = series_sum - series_term;
  assign n12897 = {1'b1, n12895};
  /* TG68K_FPU_Transcendental.vhd:1227:73  */
  assign n12898 = n12891 ? n12897 : series_term;
  /* TG68K_FPU_Transcendental.vhd:1227:73  */
  assign n12899 = n12891 ? n12896 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:1220:73  */
  assign n12900 = n12875 ? n12887 : n12898;
  /* TG68K_FPU_Transcendental.vhd:1220:73  */
  assign n12901 = n12875 ? n12888 : n12899;
  assign n12902 = {1'b1, n12871};
  /* TG68K_FPU_Transcendental.vhd:1213:73  */
  assign n12903 = n12861 ? n12902 : n12900;
  /* TG68K_FPU_Transcendental.vhd:1213:73  */
  assign n12904 = n12861 ? n12872 : n12901;
  /* TG68K_FPU_Transcendental.vhd:1238:108  */
  assign n12905 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1238:108  */
  assign n12907 = n12905 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1238:92  */
  assign n12908 = n12907[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1242:98  */
  assign n12909 = series_sum[79]; // extract
  /* TG68K_FPU_Transcendental.vhd:1243:97  */
  assign n12910 = series_sum[78:64]; // extract
  /* TG68K_FPU_Transcendental.vhd:1244:98  */
  assign n12911 = series_sum[63:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12913 = n12858 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12914 = n12858 ? result_sign : n12909;
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12915 = n12858 ? result_exp : n12910;
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12916 = n12858 ? result_mant : n12911;
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12917 = n12858 ? n12903 : series_term;
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12918 = n12858 ? n12904 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12919 = n12858 ? n12908 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:1211:65  */
  assign n12921 = n12858 ? 1'b1 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12922 = n12804 ? n12843 : n12913;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12923 = n12804 ? n12845 : n12914;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12924 = n12804 ? n12847 : n12915;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12925 = n12804 ? n12849 : n12916;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12926 = n12804 ? n12850 : n12917;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12927 = n12804 ? n12851 : n12918;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12928 = n12804 ? n12852 : n12919;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12929 = n12804 ? trans_inexact : n12921;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12930 = n12807 & n12804;
  /* TG68K_FPU_Transcendental.vhd:1182:65  */
  assign n12931 = n12804 ? n12855 : log_argument;
  /* TG68K_FPU_Transcendental.vhd:1180:57  */
  assign n12933 = operation_code == 7'b0000101;
  /* TG68K_FPU_Transcendental.vhd:1250:84  */
  assign n12934 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1250:84  */
  assign n12936 = n12934 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1258:116  */
  assign n12937 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1258:116  */
  assign n12939 = n12937 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1258:100  */
  assign n12940 = n12939[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1251:73  */
  assign n12942 = input_zero ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:1251:73  */
  assign n12944 = input_zero ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:1251:73  */
  assign n12946 = input_zero ? 15'b011111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:1251:73  */
  assign n12948 = input_zero ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:1251:73  */
  assign n12949 = input_zero ? iteration_count : n12940;
  /* TG68K_FPU_Transcendental.vhd:1260:87  */
  assign n12950 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1260:87  */
  assign n12952 = $signed(n12950) < $signed(32'b00000000000000000000000000000110);
  /* TG68K_FPU_Transcendental.vhd:1261:108  */
  assign n12953 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1261:108  */
  assign n12955 = n12953 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1261:92  */
  assign n12956 = n12955[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1265:117  */
  assign n12958 = $unsigned(input_exp) > $unsigned(15'b100000000000010);
  /* TG68K_FPU_Transcendental.vhd:1265:93  */
  assign n12959 = n12958 & input_sign;
  /* TG68K_FPU_Transcendental.vhd:1271:90  */
  assign n12960 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:1271:120  */
  assign n12962 = $unsigned(input_exp) > $unsigned(15'b100000000000010);
  /* TG68K_FPU_Transcendental.vhd:1271:96  */
  assign n12963 = n12962 & n12960;
  /* TG68K_FPU_Transcendental.vhd:1280:171  */
  assign n12964 = input_mant[63:50]; // extract
  /* TG68K_FPU_Transcendental.vhd:1280:145  */
  assign n12965 = {1'b0, n12964};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1280:143  */
  assign n12967 = 15'b011111111111111 + n12965;
  /* TG68K_FPU_Transcendental.vhd:1271:73  */
  assign n12969 = n12963 ? 15'b111111111111111 : n12967;
  /* TG68K_FPU_Transcendental.vhd:1271:73  */
  assign n12971 = n12963 ? 1'b1 : trans_overflow;
  /* TG68K_FPU_Transcendental.vhd:1265:73  */
  assign n12973 = n12959 ? 15'b000000000000000 : n12969;
  /* TG68K_FPU_Transcendental.vhd:1265:73  */
  assign n12974 = n12959 ? trans_overflow : n12971;
  /* TG68K_FPU_Transcendental.vhd:1265:73  */
  assign n12976 = n12959 ? 1'b1 : trans_underflow;
  /* TG68K_FPU_Transcendental.vhd:1260:65  */
  assign n12978 = n12952 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1260:65  */
  assign n12980 = n12952 ? result_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:1260:65  */
  assign n12981 = n12952 ? result_exp : n12973;
  /* TG68K_FPU_Transcendental.vhd:1260:65  */
  assign n12983 = n12952 ? result_mant : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1260:65  */
  assign n12984 = n12952 ? n12956 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:1260:65  */
  assign n12985 = n12952 ? trans_overflow : n12974;
  /* TG68K_FPU_Transcendental.vhd:1260:65  */
  assign n12986 = n12952 ? trans_underflow : n12976;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12987 = n12936 ? n12942 : n12978;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12988 = n12936 ? n12944 : n12980;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12989 = n12936 ? n12946 : n12981;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12990 = n12936 ? n12948 : n12983;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12991 = n12936 ? n12949 : n12984;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12992 = n12936 ? trans_overflow : n12985;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12993 = n12936 ? trans_underflow : n12986;
  /* TG68K_FPU_Transcendental.vhd:1250:65  */
  assign n12995 = n12936 ? trans_inexact : 1'b1;
  /* TG68K_FPU_Transcendental.vhd:1248:57  */
  assign n12997 = operation_code == 7'b0010001;
  /* TG68K_FPU_Transcendental.vhd:1289:84  */
  assign n12998 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1289:84  */
  assign n13000 = n12998 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1297:116  */
  assign n13001 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1297:116  */
  assign n13003 = n13001 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1297:100  */
  assign n13004 = n13003[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1290:73  */
  assign n13006 = input_zero ? 3'b111 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:1290:73  */
  assign n13008 = input_zero ? 1'b0 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:1290:73  */
  assign n13010 = input_zero ? 15'b011111111111111 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:1290:73  */
  assign n13012 = input_zero ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:1290:73  */
  assign n13013 = input_zero ? iteration_count : n13004;
  /* TG68K_FPU_Transcendental.vhd:1299:87  */
  assign n13014 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1299:87  */
  assign n13016 = $signed(n13014) < $signed(32'b00000000000000000000000000000110);
  /* TG68K_FPU_Transcendental.vhd:1300:108  */
  assign n13017 = {28'b0, iteration_count};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1300:108  */
  assign n13019 = n13017 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1300:92  */
  assign n13020 = n13019[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1304:117  */
  assign n13022 = $unsigned(input_exp) > $unsigned(15'b100000000000001);
  /* TG68K_FPU_Transcendental.vhd:1304:93  */
  assign n13023 = n13022 & input_sign;
  /* TG68K_FPU_Transcendental.vhd:1310:90  */
  assign n13024 = ~input_sign;
  /* TG68K_FPU_Transcendental.vhd:1310:120  */
  assign n13026 = $unsigned(input_exp) > $unsigned(15'b100000000000001);
  /* TG68K_FPU_Transcendental.vhd:1310:96  */
  assign n13027 = n13026 & n13024;
  /* TG68K_FPU_Transcendental.vhd:1319:183  */
  assign n13028 = input_mant[63:49]; // extract
  /* TG68K_FPU_Transcendental.vhd:1319:152  */
  assign n13030 = n13028 >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1319:143  */
  assign n13032 = 15'b011111111111111 + n13030;
  /* TG68K_FPU_Transcendental.vhd:1310:73  */
  assign n13034 = n13027 ? 15'b111111111111111 : n13032;
  /* TG68K_FPU_Transcendental.vhd:1310:73  */
  assign n13036 = n13027 ? 1'b1 : trans_overflow;
  /* TG68K_FPU_Transcendental.vhd:1304:73  */
  assign n13038 = n13023 ? 15'b000000000000000 : n13034;
  /* TG68K_FPU_Transcendental.vhd:1304:73  */
  assign n13039 = n13023 ? trans_overflow : n13036;
  /* TG68K_FPU_Transcendental.vhd:1304:73  */
  assign n13041 = n13023 ? 1'b1 : trans_underflow;
  /* TG68K_FPU_Transcendental.vhd:1299:65  */
  assign n13043 = n13016 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1299:65  */
  assign n13045 = n13016 ? result_sign : 1'b0;
  /* TG68K_FPU_Transcendental.vhd:1299:65  */
  assign n13046 = n13016 ? result_exp : n13038;
  /* TG68K_FPU_Transcendental.vhd:1299:65  */
  assign n13048 = n13016 ? result_mant : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1299:65  */
  assign n13049 = n13016 ? n13020 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:1299:65  */
  assign n13050 = n13016 ? trans_overflow : n13039;
  /* TG68K_FPU_Transcendental.vhd:1299:65  */
  assign n13051 = n13016 ? trans_underflow : n13041;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13052 = n13000 ? n13006 : n13043;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13053 = n13000 ? n13008 : n13045;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13054 = n13000 ? n13010 : n13046;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13055 = n13000 ? n13012 : n13048;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13056 = n13000 ? n13013 : n13049;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13057 = n13000 ? trans_overflow : n13050;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13058 = n13000 ? trans_underflow : n13051;
  /* TG68K_FPU_Transcendental.vhd:1289:65  */
  assign n13060 = n13000 ? trans_inexact : 1'b1;
  /* TG68K_FPU_Transcendental.vhd:1287:57  */
  assign n13062 = operation_code == 7'b0010010;
  assign n13063 = {n13062, n12997, n12933, n12801, n12671, n12533, n12482, n12462, n12262, n12095, n11946, n11810, n11677, n11539, n11509, n11479, n11376, n11361, n11349};
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13065 = n13052;
      19'b0100000000000000000: n13065 = n12987;
      19'b0010000000000000000: n13065 = n12922;
      19'b0001000000000000000: n13065 = n12789;
      19'b0000100000000000000: n13065 = n12659;
      19'b0000010000000000000: n13065 = n12524;
      19'b0000001000000000000: n13065 = n12474;
      19'b0000000100000000000: n13065 = n12448;
      19'b0000000010000000000: n13065 = n12248;
      19'b0000000001000000000: n13065 = n12082;
      19'b0000000000100000000: n13065 = n11934;
      19'b0000000000010000000: n13065 = n11797;
      19'b0000000000001000000: n13065 = n11664;
      19'b0000000000000100000: n13065 = n11532;
      19'b0000000000000010000: n13065 = n11502;
      19'b0000000000000001000: n13065 = n11469;
      19'b0000000000000000100: n13065 = n11366;
      19'b0000000000000000010: n13065 = n11354;
      19'b0000000000000000001: n13065 = n11337;
      default: n13065 = 3'b111;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13066 = cordic_iteration;
      19'b0100000000000000000: n13066 = cordic_iteration;
      19'b0010000000000000000: n13066 = cordic_iteration;
      19'b0001000000000000000: n13066 = cordic_iteration;
      19'b0000100000000000000: n13066 = cordic_iteration;
      19'b0000010000000000000: n13066 = cordic_iteration;
      19'b0000001000000000000: n13066 = n12475;
      19'b0000000100000000000: n13066 = cordic_iteration;
      19'b0000000010000000000: n13066 = cordic_iteration;
      19'b0000000001000000000: n13066 = cordic_iteration;
      19'b0000000000100000000: n13066 = cordic_iteration;
      19'b0000000000010000000: n13066 = cordic_iteration;
      19'b0000000000001000000: n13066 = cordic_iteration;
      19'b0000000000000100000: n13066 = cordic_iteration;
      19'b0000000000000010000: n13066 = cordic_iteration;
      19'b0000000000000001000: n13066 = cordic_iteration;
      19'b0000000000000000100: n13066 = n11368;
      19'b0000000000000000010: n13066 = n11356;
      19'b0000000000000000001: n13066 = cordic_iteration;
      default: n13066 = cordic_iteration;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13068 = n13053;
      19'b0100000000000000000: n13068 = n12988;
      19'b0010000000000000000: n13068 = n12923;
      19'b0001000000000000000: n13068 = n12790;
      19'b0000100000000000000: n13068 = n12660;
      19'b0000010000000000000: n13068 = n12525;
      19'b0000001000000000000: n13068 = n12476;
      19'b0000000100000000000: n13068 = n12449;
      19'b0000000010000000000: n13068 = n12249;
      19'b0000000001000000000: n13068 = n12083;
      19'b0000000000100000000: n13068 = n11935;
      19'b0000000000010000000: n13068 = n11798;
      19'b0000000000001000000: n13068 = n11665;
      19'b0000000000000100000: n13068 = n11534;
      19'b0000000000000010000: n13068 = n11504;
      19'b0000000000000001000: n13068 = n11470;
      19'b0000000000000000100: n13068 = n11370;
      19'b0000000000000000010: n13068 = n11357;
      19'b0000000000000000001: n13068 = n11338;
      default: n13068 = 1'b0;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13070 = n13054;
      19'b0100000000000000000: n13070 = n12989;
      19'b0010000000000000000: n13070 = n12924;
      19'b0001000000000000000: n13070 = n12791;
      19'b0000100000000000000: n13070 = n12661;
      19'b0000010000000000000: n13070 = n12526;
      19'b0000001000000000000: n13070 = n12478;
      19'b0000000100000000000: n13070 = n12450;
      19'b0000000010000000000: n13070 = n12250;
      19'b0000000001000000000: n13070 = n12084;
      19'b0000000000100000000: n13070 = n11936;
      19'b0000000000010000000: n13070 = n11799;
      19'b0000000000001000000: n13070 = n11666;
      19'b0000000000000100000: n13070 = n11535;
      19'b0000000000000010000: n13070 = n11505;
      19'b0000000000000001000: n13070 = n11471;
      19'b0000000000000000100: n13070 = n11372;
      19'b0000000000000000010: n13070 = n11358;
      19'b0000000000000000001: n13070 = n11339;
      default: n13070 = 15'b111111111111111;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13072 = n13055;
      19'b0100000000000000000: n13072 = n12990;
      19'b0010000000000000000: n13072 = n12925;
      19'b0001000000000000000: n13072 = n12792;
      19'b0000100000000000000: n13072 = n12662;
      19'b0000010000000000000: n13072 = n12527;
      19'b0000001000000000000: n13072 = n12480;
      19'b0000000100000000000: n13072 = n12451;
      19'b0000000010000000000: n13072 = n12251;
      19'b0000000001000000000: n13072 = n12085;
      19'b0000000000100000000: n13072 = n11937;
      19'b0000000000010000000: n13072 = n11800;
      19'b0000000000001000000: n13072 = n11667;
      19'b0000000000000100000: n13072 = n11536;
      19'b0000000000000010000: n13072 = n11506;
      19'b0000000000000001000: n13072 = n11472;
      19'b0000000000000000100: n13072 = n11374;
      19'b0000000000000000010: n13072 = n11359;
      19'b0000000000000000001: n13072 = n11340;
      default: n13072 = 64'b1100000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13073 = series_term;
      19'b0100000000000000000: n13073 = series_term;
      19'b0010000000000000000: n13073 = n12926;
      19'b0001000000000000000: n13073 = n12793;
      19'b0000100000000000000: n13073 = n12663;
      19'b0000010000000000000: n13073 = series_term;
      19'b0000001000000000000: n13073 = series_term;
      19'b0000000100000000000: n13073 = series_term;
      19'b0000000010000000000: n13073 = series_term;
      19'b0000000001000000000: n13073 = series_term;
      19'b0000000000100000000: n13073 = series_term;
      19'b0000000000010000000: n13073 = series_term;
      19'b0000000000001000000: n13073 = series_term;
      19'b0000000000000100000: n13073 = series_term;
      19'b0000000000000010000: n13073 = series_term;
      19'b0000000000000001000: n13073 = n11473;
      19'b0000000000000000100: n13073 = series_term;
      19'b0000000000000000010: n13073 = series_term;
      19'b0000000000000000001: n13073 = series_term;
      default: n13073 = series_term;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13074 = series_sum;
      19'b0100000000000000000: n13074 = series_sum;
      19'b0010000000000000000: n13074 = n12927;
      19'b0001000000000000000: n13074 = n12794;
      19'b0000100000000000000: n13074 = n12664;
      19'b0000010000000000000: n13074 = series_sum;
      19'b0000001000000000000: n13074 = series_sum;
      19'b0000000100000000000: n13074 = n12452;
      19'b0000000010000000000: n13074 = n12252;
      19'b0000000001000000000: n13074 = n12086;
      19'b0000000000100000000: n13074 = n11938;
      19'b0000000000010000000: n13074 = n11801;
      19'b0000000000001000000: n13074 = n11668;
      19'b0000000000000100000: n13074 = series_sum;
      19'b0000000000000010000: n13074 = series_sum;
      19'b0000000000000001000: n13074 = n11474;
      19'b0000000000000000100: n13074 = series_sum;
      19'b0000000000000000010: n13074 = series_sum;
      19'b0000000000000000001: n13074 = series_sum;
      default: n13074 = series_sum;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13075 = n13056;
      19'b0100000000000000000: n13075 = n12991;
      19'b0010000000000000000: n13075 = n12928;
      19'b0001000000000000000: n13075 = n12795;
      19'b0000100000000000000: n13075 = n12665;
      19'b0000010000000000000: n13075 = n12528;
      19'b0000001000000000000: n13075 = iteration_count;
      19'b0000000100000000000: n13075 = n12453;
      19'b0000000010000000000: n13075 = n12253;
      19'b0000000001000000000: n13075 = n12087;
      19'b0000000000100000000: n13075 = n11939;
      19'b0000000000010000000: n13075 = n11802;
      19'b0000000000001000000: n13075 = n11669;
      19'b0000000000000100000: n13075 = n11537;
      19'b0000000000000010000: n13075 = n11507;
      19'b0000000000000001000: n13075 = n11475;
      19'b0000000000000000100: n13075 = iteration_count;
      19'b0000000000000000010: n13075 = iteration_count;
      19'b0000000000000000001: n13075 = n11341;
      default: n13075 = iteration_count;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13076 = n13057;
      19'b0100000000000000000: n13076 = n12992;
      19'b0010000000000000000: n13076 = trans_overflow;
      19'b0001000000000000000: n13076 = n12796;
      19'b0000100000000000000: n13076 = n12666;
      19'b0000010000000000000: n13076 = trans_overflow;
      19'b0000001000000000000: n13076 = trans_overflow;
      19'b0000000100000000000: n13076 = trans_overflow;
      19'b0000000010000000000: n13076 = trans_overflow;
      19'b0000000001000000000: n13076 = trans_overflow;
      19'b0000000000100000000: n13076 = trans_overflow;
      19'b0000000000010000000: n13076 = trans_overflow;
      19'b0000000000001000000: n13076 = trans_overflow;
      19'b0000000000000100000: n13076 = trans_overflow;
      19'b0000000000000010000: n13076 = trans_overflow;
      19'b0000000000000001000: n13076 = trans_overflow;
      19'b0000000000000000100: n13076 = trans_overflow;
      19'b0000000000000000010: n13076 = trans_overflow;
      19'b0000000000000000001: n13076 = trans_overflow;
      default: n13076 = trans_overflow;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13077 = n13058;
      19'b0100000000000000000: n13077 = n12993;
      19'b0010000000000000000: n13077 = trans_underflow;
      19'b0001000000000000000: n13077 = n12797;
      19'b0000100000000000000: n13077 = n12667;
      19'b0000010000000000000: n13077 = trans_underflow;
      19'b0000001000000000000: n13077 = trans_underflow;
      19'b0000000100000000000: n13077 = trans_underflow;
      19'b0000000010000000000: n13077 = trans_underflow;
      19'b0000000001000000000: n13077 = trans_underflow;
      19'b0000000000100000000: n13077 = trans_underflow;
      19'b0000000000010000000: n13077 = trans_underflow;
      19'b0000000000001000000: n13077 = trans_underflow;
      19'b0000000000000100000: n13077 = trans_underflow;
      19'b0000000000000010000: n13077 = trans_underflow;
      19'b0000000000000001000: n13077 = trans_underflow;
      19'b0000000000000000100: n13077 = trans_underflow;
      19'b0000000000000000010: n13077 = trans_underflow;
      19'b0000000000000000001: n13077 = trans_underflow;
      default: n13077 = trans_underflow;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13080 = n13060;
      19'b0100000000000000000: n13080 = n12995;
      19'b0010000000000000000: n13080 = n12929;
      19'b0001000000000000000: n13080 = n12798;
      19'b0000100000000000000: n13080 = n12668;
      19'b0000010000000000000: n13080 = n12530;
      19'b0000001000000000000: n13080 = trans_inexact;
      19'b0000000100000000000: n13080 = n12454;
      19'b0000000010000000000: n13080 = n12254;
      19'b0000000001000000000: n13080 = n12088;
      19'b0000000000100000000: n13080 = n11940;
      19'b0000000000010000000: n13080 = n11803;
      19'b0000000000001000000: n13080 = n11670;
      19'b0000000000000100000: n13080 = 1'b1;
      19'b0000000000000010000: n13080 = 1'b1;
      19'b0000000000000001000: n13080 = n11476;
      19'b0000000000000000100: n13080 = trans_inexact;
      19'b0000000000000000010: n13080 = trans_inexact;
      19'b0000000000000000001: n13080 = n11342;
      default: n13080 = trans_inexact;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13082 = trans_invalid;
      19'b0100000000000000000: n13082 = trans_invalid;
      19'b0010000000000000000: n13082 = n12854;
      19'b0001000000000000000: n13082 = trans_invalid;
      19'b0000100000000000000: n13082 = trans_invalid;
      19'b0000010000000000000: n13082 = n12510;
      19'b0000001000000000000: n13082 = trans_invalid;
      19'b0000000100000000000: n13082 = n12335;
      19'b0000000010000000000: n13082 = n12146;
      19'b0000000001000000000: n13082 = trans_invalid;
      19'b0000000000100000000: n13082 = trans_invalid;
      19'b0000000000010000000: n13082 = trans_invalid;
      19'b0000000000001000000: n13082 = trans_invalid;
      19'b0000000000000100000: n13082 = trans_invalid;
      19'b0000000000000010000: n13082 = trans_invalid;
      19'b0000000000000001000: n13082 = trans_invalid;
      19'b0000000000000000100: n13082 = trans_invalid;
      19'b0000000000000000010: n13082 = trans_invalid;
      19'b0000000000000000001: n13082 = trans_invalid;
      default: n13082 = 1'b1;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13083 = exp_argument;
      19'b0100000000000000000: n13083 = exp_argument;
      19'b0010000000000000000: n13083 = exp_argument;
      19'b0001000000000000000: n13083 = n12799;
      19'b0000100000000000000: n13083 = n12669;
      19'b0000010000000000000: n13083 = exp_argument;
      19'b0000001000000000000: n13083 = exp_argument;
      19'b0000000100000000000: n13083 = exp_argument;
      19'b0000000010000000000: n13083 = exp_argument;
      19'b0000000001000000000: n13083 = exp_argument;
      19'b0000000000100000000: n13083 = exp_argument;
      19'b0000000000010000000: n13083 = exp_argument;
      19'b0000000000001000000: n13083 = exp_argument;
      19'b0000000000000100000: n13083 = exp_argument;
      19'b0000000000000010000: n13083 = exp_argument;
      19'b0000000000000001000: n13083 = exp_argument;
      19'b0000000000000000100: n13083 = exp_argument;
      19'b0000000000000000010: n13083 = exp_argument;
      19'b0000000000000000001: n13083 = exp_argument;
      default: n13083 = exp_argument;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13084 = log_argument;
      19'b0100000000000000000: n13084 = log_argument;
      19'b0010000000000000000: n13084 = n12931;
      19'b0001000000000000000: n13084 = log_argument;
      19'b0000100000000000000: n13084 = log_argument;
      19'b0000010000000000000: n13084 = log_argument;
      19'b0000001000000000000: n13084 = log_argument;
      19'b0000000100000000000: n13084 = log_argument;
      19'b0000000010000000000: n13084 = log_argument;
      19'b0000000001000000000: n13084 = log_argument;
      19'b0000000000100000000: n13084 = log_argument;
      19'b0000000000010000000: n13084 = log_argument;
      19'b0000000000001000000: n13084 = log_argument;
      19'b0000000000000100000: n13084 = log_argument;
      19'b0000000000000010000: n13084 = log_argument;
      19'b0000000000000001000: n13084 = n11477;
      19'b0000000000000000100: n13084 = log_argument;
      19'b0000000000000000010: n13084 = log_argument;
      19'b0000000000000000001: n13084 = log_argument;
      default: n13084 = log_argument;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13085 = x_squared;
      19'b0100000000000000000: n13085 = x_squared;
      19'b0010000000000000000: n13085 = x_squared;
      19'b0001000000000000000: n13085 = x_squared;
      19'b0000100000000000000: n13085 = x_squared;
      19'b0000010000000000000: n13085 = x_squared;
      19'b0000001000000000000: n13085 = x_squared;
      19'b0000000100000000000: n13085 = n12456;
      19'b0000000010000000000: n13085 = n12256;
      19'b0000000001000000000: n13085 = n12089;
      19'b0000000000100000000: n13085 = n11941;
      19'b0000000000010000000: n13085 = n11804;
      19'b0000000000001000000: n13085 = n11671;
      19'b0000000000000100000: n13085 = x_squared;
      19'b0000000000000010000: n13085 = x_squared;
      19'b0000000000000001000: n13085 = x_squared;
      19'b0000000000000000100: n13085 = x_squared;
      19'b0000000000000000010: n13085 = x_squared;
      19'b0000000000000000001: n13085 = x_squared;
      default: n13085 = x_squared;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13086 = x_cubed;
      19'b0100000000000000000: n13086 = x_cubed;
      19'b0010000000000000000: n13086 = x_cubed;
      19'b0001000000000000000: n13086 = x_cubed;
      19'b0000100000000000000: n13086 = x_cubed;
      19'b0000010000000000000: n13086 = x_cubed;
      19'b0000001000000000000: n13086 = x_cubed;
      19'b0000000100000000000: n13086 = n12457;
      19'b0000000010000000000: n13086 = n12257;
      19'b0000000001000000000: n13086 = n12090;
      19'b0000000000100000000: n13086 = n11942;
      19'b0000000000010000000: n13086 = n11805;
      19'b0000000000001000000: n13086 = n11672;
      19'b0000000000000100000: n13086 = x_cubed;
      19'b0000000000000010000: n13086 = x_cubed;
      19'b0000000000000001000: n13086 = x_cubed;
      19'b0000000000000000100: n13086 = x_cubed;
      19'b0000000000000000010: n13086 = x_cubed;
      19'b0000000000000000001: n13086 = x_cubed;
      default: n13086 = x_cubed;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13087 = x_fifth;
      19'b0100000000000000000: n13087 = x_fifth;
      19'b0010000000000000000: n13087 = x_fifth;
      19'b0001000000000000000: n13087 = x_fifth;
      19'b0000100000000000000: n13087 = x_fifth;
      19'b0000010000000000000: n13087 = x_fifth;
      19'b0000001000000000000: n13087 = x_fifth;
      19'b0000000100000000000: n13087 = n12458;
      19'b0000000010000000000: n13087 = n12258;
      19'b0000000001000000000: n13087 = n12091;
      19'b0000000000100000000: n13087 = n11943;
      19'b0000000000010000000: n13087 = n11806;
      19'b0000000000001000000: n13087 = n11673;
      19'b0000000000000100000: n13087 = x_fifth;
      19'b0000000000000010000: n13087 = x_fifth;
      19'b0000000000000001000: n13087 = x_fifth;
      19'b0000000000000000100: n13087 = x_fifth;
      19'b0000000000000000010: n13087 = x_fifth;
      19'b0000000000000000001: n13087 = x_fifth;
      default: n13087 = x_fifth;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13088 = x3_div6;
      19'b0100000000000000000: n13088 = x3_div6;
      19'b0010000000000000000: n13088 = x3_div6;
      19'b0001000000000000000: n13088 = x3_div6;
      19'b0000100000000000000: n13088 = x3_div6;
      19'b0000010000000000000: n13088 = x3_div6;
      19'b0000001000000000000: n13088 = x3_div6;
      19'b0000000100000000000: n13088 = n12459;
      19'b0000000010000000000: n13088 = n12259;
      19'b0000000001000000000: n13088 = n12092;
      19'b0000000000100000000: n13088 = x3_div6;
      19'b0000000000010000000: n13088 = n11807;
      19'b0000000000001000000: n13088 = n11674;
      19'b0000000000000100000: n13088 = x3_div6;
      19'b0000000000000010000: n13088 = x3_div6;
      19'b0000000000000001000: n13088 = x3_div6;
      19'b0000000000000000100: n13088 = x3_div6;
      19'b0000000000000000010: n13088 = x3_div6;
      19'b0000000000000000001: n13088 = x3_div6;
      default: n13088 = x3_div6;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13089 = x5_div120;
      19'b0100000000000000000: n13089 = x5_div120;
      19'b0010000000000000000: n13089 = x5_div120;
      19'b0001000000000000000: n13089 = x5_div120;
      19'b0000100000000000000: n13089 = x5_div120;
      19'b0000010000000000000: n13089 = x5_div120;
      19'b0000001000000000000: n13089 = x5_div120;
      19'b0000000100000000000: n13089 = n12460;
      19'b0000000010000000000: n13089 = n12260;
      19'b0000000001000000000: n13089 = n12093;
      19'b0000000000100000000: n13089 = n11944;
      19'b0000000000010000000: n13089 = n11808;
      19'b0000000000001000000: n13089 = n11675;
      19'b0000000000000100000: n13089 = x5_div120;
      19'b0000000000000010000: n13089 = x5_div120;
      19'b0000000000000001000: n13089 = x5_div120;
      19'b0000000000000000100: n13089 = x5_div120;
      19'b0000000000000000010: n13089 = x5_div120;
      19'b0000000000000000001: n13089 = x5_div120;
      default: n13089 = x5_div120;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13090 = x_n;
      19'b0100000000000000000: n13090 = x_n;
      19'b0010000000000000000: n13090 = x_n;
      19'b0001000000000000000: n13090 = x_n;
      19'b0000100000000000000: n13090 = x_n;
      19'b0000010000000000000: n13090 = x_n;
      19'b0000001000000000000: n13090 = x_n;
      19'b0000000100000000000: n13090 = x_n;
      19'b0000000010000000000: n13090 = x_n;
      19'b0000000001000000000: n13090 = x_n;
      19'b0000000000100000000: n13090 = x_n;
      19'b0000000000010000000: n13090 = x_n;
      19'b0000000000001000000: n13090 = x_n;
      19'b0000000000000100000: n13090 = x_n;
      19'b0000000000000010000: n13090 = x_n;
      19'b0000000000000001000: n13090 = x_n;
      19'b0000000000000000100: n13090 = x_n;
      19'b0000000000000000010: n13090 = x_n;
      19'b0000000000000000001: n13090 = n11344;
      default: n13090 = x_n;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13091 = a_div_x_n;
      19'b0100000000000000000: n13091 = a_div_x_n;
      19'b0010000000000000000: n13091 = a_div_x_n;
      19'b0001000000000000000: n13091 = a_div_x_n;
      19'b0000100000000000000: n13091 = a_div_x_n;
      19'b0000010000000000000: n13091 = a_div_x_n;
      19'b0000001000000000000: n13091 = a_div_x_n;
      19'b0000000100000000000: n13091 = a_div_x_n;
      19'b0000000010000000000: n13091 = a_div_x_n;
      19'b0000000001000000000: n13091 = a_div_x_n;
      19'b0000000000100000000: n13091 = a_div_x_n;
      19'b0000000000010000000: n13091 = a_div_x_n;
      19'b0000000000001000000: n13091 = a_div_x_n;
      19'b0000000000000100000: n13091 = a_div_x_n;
      19'b0000000000000010000: n13091 = a_div_x_n;
      19'b0000000000000001000: n13091 = a_div_x_n;
      19'b0000000000000000100: n13091 = a_div_x_n;
      19'b0000000000000000010: n13091 = a_div_x_n;
      19'b0000000000000000001: n13091 = n11345;
      default: n13091 = a_div_x_n;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13092 = x_next;
      19'b0100000000000000000: n13092 = x_next;
      19'b0010000000000000000: n13092 = x_next;
      19'b0001000000000000000: n13092 = x_next;
      19'b0000100000000000000: n13092 = x_next;
      19'b0000010000000000000: n13092 = x_next;
      19'b0000001000000000000: n13092 = x_next;
      19'b0000000100000000000: n13092 = x_next;
      19'b0000000010000000000: n13092 = x_next;
      19'b0000000001000000000: n13092 = x_next;
      19'b0000000000100000000: n13092 = x_next;
      19'b0000000000010000000: n13092 = x_next;
      19'b0000000000001000000: n13092 = x_next;
      19'b0000000000000100000: n13092 = x_next;
      19'b0000000000000010000: n13092 = x_next;
      19'b0000000000000001000: n13092 = x_next;
      19'b0000000000000000100: n13092 = x_next;
      19'b0000000000000000010: n13092 = x_next;
      19'b0000000000000000001: n13092 = n11346;
      default: n13092 = x_next;
    endcase
  /* TG68K_FPU_Transcendental.vhd:356:49  */
  always @*
    case (n13063)
      19'b1000000000000000000: n13093 = final_mant;
      19'b0100000000000000000: n13093 = final_mant;
      19'b0010000000000000000: n13093 = final_mant;
      19'b0001000000000000000: n13093 = final_mant;
      19'b0000100000000000000: n13093 = final_mant;
      19'b0000010000000000000: n13093 = final_mant;
      19'b0000001000000000000: n13093 = final_mant;
      19'b0000000100000000000: n13093 = final_mant;
      19'b0000000010000000000: n13093 = final_mant;
      19'b0000000001000000000: n13093 = final_mant;
      19'b0000000000100000000: n13093 = final_mant;
      19'b0000000000010000000: n13093 = final_mant;
      19'b0000000000001000000: n13093 = final_mant;
      19'b0000000000000100000: n13093 = final_mant;
      19'b0000000000000010000: n13093 = final_mant;
      19'b0000000000000001000: n13093 = final_mant;
      19'b0000000000000000100: n13093 = final_mant;
      19'b0000000000000000010: n13093 = final_mant;
      19'b0000000000000000001: n13093 = n11347;
      default: n13093 = final_mant;
    endcase
  /* TG68K_FPU_Transcendental.vhd:354:41  */
  assign n13095 = trans_state == 3'b011;
  /* TG68K_FPU_Transcendental.vhd:1335:41  */
  assign n13097 = trans_state == 3'b100;
  /* TG68K_FPU_Transcendental.vhd:1341:69  */
  assign n13098 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1341:69  */
  assign n13100 = n13098 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1350:118  */
  assign n13101 = input_mant[63:34]; // extract
  /* TG68K_FPU_Transcendental.vhd:1350:92  */
  assign n13102 = {34'b0, n13101};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1352:110  */
  assign n13103 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1352:110  */
  assign n13105 = n13103 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1352:93  */
  assign n13106 = n13105[4:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1344:65  */
  assign n13108 = operation_code == 7'b0001110;
  /* TG68K_FPU_Transcendental.vhd:1344:78  */
  assign n13110 = operation_code == 7'b0011101;
  /* TG68K_FPU_Transcendental.vhd:1344:78  */
  assign n13111 = n13108 | n13110;
  /* TG68K_FPU_Transcendental.vhd:1355:118  */
  assign n13112 = input_mant[63:34]; // extract
  /* TG68K_FPU_Transcendental.vhd:1355:92  */
  assign n13113 = {34'b0, n13112};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1356:115  */
  assign n13114 = operand[39:10]; // extract
  /* TG68K_FPU_Transcendental.vhd:1356:92  */
  assign n13115 = {34'b0, n13114};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1359:110  */
  assign n13116 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1359:110  */
  assign n13118 = n13116 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1359:93  */
  assign n13119 = n13118[4:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1353:65  */
  assign n13121 = operation_code == 7'b0001010;
  assign n13122 = {n13121, n13111};
  /* TG68K_FPU_Transcendental.vhd:1343:57  */
  always @*
    case (n13122)
      2'b10: n13124 = trans_state;
      2'b01: n13124 = trans_state;
      default: n13124 = 3'b110;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1343:57  */
  always @*
    case (n13122)
      2'b10: n13126 = n13113;
      2'b01: n13126 = 64'b0000000000000000000000000000000001101010000010011110011001100111;
      default: n13126 = cordic_x;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1343:57  */
  always @*
    case (n13122)
      2'b10: n13128 = n13115;
      2'b01: n13128 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      default: n13128 = cordic_y;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1343:57  */
  always @*
    case (n13122)
      2'b10: n13130 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      2'b01: n13130 = n13102;
      default: n13130 = cordic_z;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1343:57  */
  always @*
    case (n13122)
      2'b10: n13131 = n13119;
      2'b01: n13131 = n13106;
      default: n13131 = cordic_iteration;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1343:57  */
  always @*
    case (n13122)
      2'b10: n13134 = 1'b1;
      2'b01: n13134 = 1'b0;
      default: n13134 = cordic_mode;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1364:72  */
  assign n13135 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1364:72  */
  assign n13137 = $signed(n13135) <= $signed(32'b00000000000000000000000000001111);
  /* TG68K_FPU_Transcendental.vhd:1367:114  */
  assign n13138 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1367:114  */
  assign n13140 = n13138 - 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1367:97  */
  assign n13141 = n13140[30:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1367:75  */
  assign n13142 = $signed(cordic_x) >>> n13141;
  /* TG68K_FPU_Transcendental.vhd:1368:114  */
  assign n13143 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1368:114  */
  assign n13145 = n13143 - 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1368:97  */
  assign n13146 = n13145[30:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1368:75  */
  assign n13147 = $signed(cordic_y) >>> n13146;
  /* TG68K_FPU_Transcendental.vhd:1369:118  */
  assign n13148 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1369:118  */
  assign n13150 = n13148 - 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1369:118  */
  assign n13151 = n13150[3:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1371:72  */
  assign n13157 = ~cordic_mode;
  /* TG68K_FPU_Transcendental.vhd:1373:77  */
  assign n13159 = $signed(cordic_z) >= $signed(64'b0000000000000000000000000000000000000000000000000000000000000000);
  /* TG68K_FPU_Transcendental.vhd:1375:94  */
  assign n13160 = cordic_x - cordic_shift_y;
  /* TG68K_FPU_Transcendental.vhd:1376:94  */
  assign n13161 = cordic_y + cordic_shift_x;
  /* TG68K_FPU_Transcendental.vhd:1377:94  */
  assign n13162 = cordic_z - cordic_atan_val;
  /* TG68K_FPU_Transcendental.vhd:1380:94  */
  assign n13163 = cordic_x + cordic_shift_y;
  /* TG68K_FPU_Transcendental.vhd:1381:94  */
  assign n13164 = cordic_y - cordic_shift_x;
  /* TG68K_FPU_Transcendental.vhd:1382:94  */
  assign n13165 = cordic_z + cordic_atan_val;
  /* TG68K_FPU_Transcendental.vhd:1373:65  */
  assign n13166 = n13159 ? n13160 : n13163;
  /* TG68K_FPU_Transcendental.vhd:1373:65  */
  assign n13167 = n13159 ? n13161 : n13164;
  /* TG68K_FPU_Transcendental.vhd:1373:65  */
  assign n13168 = n13159 ? n13162 : n13165;
  /* TG68K_FPU_Transcendental.vhd:1386:77  */
  assign n13170 = $signed(cordic_y) >= $signed(64'b0000000000000000000000000000000000000000000000000000000000000000);
  /* TG68K_FPU_Transcendental.vhd:1387:94  */
  assign n13171 = cordic_x + cordic_shift_y;
  /* TG68K_FPU_Transcendental.vhd:1388:94  */
  assign n13172 = cordic_y - cordic_shift_x;
  /* TG68K_FPU_Transcendental.vhd:1389:94  */
  assign n13173 = cordic_z + cordic_atan_val;
  /* TG68K_FPU_Transcendental.vhd:1391:94  */
  assign n13174 = cordic_x - cordic_shift_y;
  /* TG68K_FPU_Transcendental.vhd:1392:94  */
  assign n13175 = cordic_y + cordic_shift_x;
  /* TG68K_FPU_Transcendental.vhd:1393:94  */
  assign n13176 = cordic_z - cordic_atan_val;
  /* TG68K_FPU_Transcendental.vhd:1386:65  */
  assign n13177 = n13170 ? n13171 : n13174;
  /* TG68K_FPU_Transcendental.vhd:1386:65  */
  assign n13178 = n13170 ? n13172 : n13175;
  /* TG68K_FPU_Transcendental.vhd:1386:65  */
  assign n13179 = n13170 ? n13173 : n13176;
  /* TG68K_FPU_Transcendental.vhd:1371:57  */
  assign n13180 = n13157 ? n13166 : n13177;
  /* TG68K_FPU_Transcendental.vhd:1371:57  */
  assign n13181 = n13157 ? n13167 : n13178;
  /* TG68K_FPU_Transcendental.vhd:1371:57  */
  assign n13182 = n13157 ? n13168 : n13179;
  /* TG68K_FPU_Transcendental.vhd:1397:94  */
  assign n13183 = {27'b0, cordic_iteration};  //  uext
  /* TG68K_FPU_Transcendental.vhd:1397:94  */
  assign n13185 = n13183 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU_Transcendental.vhd:1397:77  */
  assign n13186 = n13185[4:0];  // trunc
  /* TG68K_FPU_Transcendental.vhd:1405:121  */
  assign n13187 = $signed(cordic_y) >= 0 ? cordic_y : -cordic_y;
  /* TG68K_FPU_Transcendental.vhd:1401:65  */
  assign n13189 = operation_code == 7'b0001110;
  /* TG68K_FPU_Transcendental.vhd:1410:121  */
  assign n13190 = $signed(cordic_x) >= 0 ? cordic_x : -cordic_x;
  /* TG68K_FPU_Transcendental.vhd:1406:65  */
  assign n13192 = operation_code == 7'b0011101;
  /* TG68K_FPU_Transcendental.vhd:1413:96  */
  assign n13193 = cordic_z[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:1415:121  */
  assign n13194 = $signed(cordic_z) >= 0 ? cordic_z : -cordic_z;
  /* TG68K_FPU_Transcendental.vhd:1411:65  */
  assign n13196 = operation_code == 7'b0001010;
  assign n13197 = {n13196, n13192, n13189};
  /* TG68K_FPU_Transcendental.vhd:1400:57  */
  always @*
    case (n13197)
      3'b100: n13201 = n13193;
      3'b010: n13201 = 1'b0;
      3'b001: n13201 = input_sign;
      default: n13201 = result_sign;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1400:57  */
  always @*
    case (n13197)
      3'b100: n13205 = 15'b011111111111111;
      3'b010: n13205 = 15'b011111111111110;
      3'b001: n13205 = 15'b011111111111110;
      default: n13205 = result_exp;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1400:57  */
  always @*
    case (n13197)
      3'b100: n13206 = n13194;
      3'b010: n13206 = n13190;
      3'b001: n13206 = n13187;
      default: n13206 = result_mant;
    endcase
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13208 = n13137 ? trans_state : 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13209 = n13137 ? n13180 : cordic_x;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13210 = n13137 ? n13181 : cordic_y;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13211 = n13137 ? n13182 : cordic_z;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13212 = n13137 ? n13186 : cordic_iteration;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13213 = n13137 ? result_sign : n13201;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13214 = n13137 ? result_exp : n13205;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13215 = n13137 ? result_mant : n13206;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13216 = n13137 ? n13142 : cordic_shift_x;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13217 = n13137 ? n13147 : cordic_shift_y;
  /* TG68K_FPU_Transcendental.vhd:1364:49  */
  assign n13218 = n13137 ? n13645 : cordic_atan_val;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13219 = n13100 ? n13124 : n13208;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13220 = n13100 ? n13126 : n13209;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13221 = n13100 ? n13128 : n13210;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13222 = n13100 ? n13130 : n13211;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13223 = n13100 ? n13131 : n13212;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13224 = n13100 ? n13134 : cordic_mode;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13225 = n13100 ? result_sign : n13213;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13226 = n13100 ? result_exp : n13214;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13227 = n13100 ? result_mant : n13215;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13228 = n13100 ? cordic_shift_x : n13216;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13229 = n13100 ? cordic_shift_y : n13217;
  /* TG68K_FPU_Transcendental.vhd:1341:49  */
  assign n13230 = n13100 ? cordic_atan_val : n13218;
  /* TG68K_FPU_Transcendental.vhd:1339:41  */
  assign n13232 = trans_state == 3'b101;
  /* TG68K_FPU_Transcendental.vhd:1425:63  */
  assign n13234 = result_exp == 15'b000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1425:99  */
  assign n13236 = result_mant != 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1425:83  */
  assign n13237 = n13236 & n13234;
  /* TG68K_FPU_Transcendental.vhd:1427:71  */
  assign n13238 = result_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:1427:76  */
  assign n13239 = ~n13238;
  /* TG68K_FPU_Transcendental.vhd:1429:79  */
  assign n13240 = result_mant[62]; // extract
  /* TG68K_FPU_Transcendental.vhd:1430:99  */
  assign n13241 = result_mant[62:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1430:113  */
  assign n13243 = {n13241, 1'b0};
  /* TG68K_FPU_Transcendental.vhd:1432:82  */
  assign n13244 = result_mant[61]; // extract
  /* TG68K_FPU_Transcendental.vhd:1433:99  */
  assign n13245 = result_mant[61:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1433:113  */
  assign n13247 = {n13245, 2'b00};
  /* TG68K_FPU_Transcendental.vhd:1437:99  */
  assign n13248 = result_mant[59:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1437:113  */
  assign n13250 = {n13248, 4'b0000};
  /* TG68K_FPU_Transcendental.vhd:1432:65  */
  assign n13253 = n13244 ? 15'b000000000000010 : 15'b000000000000100;
  /* TG68K_FPU_Transcendental.vhd:1432:65  */
  assign n13254 = n13244 ? n13247 : n13250;
  /* TG68K_FPU_Transcendental.vhd:1429:65  */
  assign n13256 = n13240 ? 15'b000000000000001 : n13253;
  /* TG68K_FPU_Transcendental.vhd:1429:65  */
  assign n13257 = n13240 ? n13243 : n13254;
  /* TG68K_FPU_Transcendental.vhd:1425:49  */
  assign n13258 = n13286 ? n13256 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:1427:57  */
  assign n13259 = n13239 ? n13257 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:1441:66  */
  assign n13261 = result_exp == 15'b111111111111111;
  /* TG68K_FPU_Transcendental.vhd:1443:71  */
  assign n13262 = result_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:1443:97  */
  assign n13263 = result_mant[62:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1443:111  */
  assign n13265 = n13263 == 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_Transcendental.vhd:1443:82  */
  assign n13266 = n13265 & n13262;
  assign n13268 = result_mant[62]; // extract
  /* TG68K_FPU_Transcendental.vhd:1443:57  */
  assign n13269 = n13266 ? n13268 : 1'b1;
  /* TG68K_FPU_Transcendental.vhd:1450:76  */
  assign n13271 = $unsigned(result_exp) > $unsigned(15'b000000000000000);
  /* TG68K_FPU_Transcendental.vhd:1450:105  */
  assign n13273 = $unsigned(result_exp) < $unsigned(15'b111111111111111);
  /* TG68K_FPU_Transcendental.vhd:1450:80  */
  assign n13274 = n13273 & n13271;
  /* TG68K_FPU_Transcendental.vhd:1452:71  */
  assign n13275 = result_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:1452:76  */
  assign n13276 = ~n13275;
  assign n13278 = result_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:1450:49  */
  assign n13279 = n13281 ? 1'b1 : n13278;
  /* TG68K_FPU_Transcendental.vhd:1450:49  */
  assign n13281 = n13276 & n13274;
  assign n13282 = result_mant[62]; // extract
  /* TG68K_FPU_Transcendental.vhd:1441:49  */
  assign n13283 = n13261 ? n13269 : n13282;
  assign n13284 = result_mant[63]; // extract
  /* TG68K_FPU_Transcendental.vhd:1441:49  */
  assign n13285 = n13261 ? n13284 : n13279;
  /* TG68K_FPU_Transcendental.vhd:1425:49  */
  assign n13286 = n13239 & n13237;
  assign n13287 = {n13285, n13283};
  assign n13288 = n13259[61:0]; // extract
  assign n13289 = result_mant[61:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:1425:49  */
  assign n13290 = n13237 ? n13288 : n13289;
  assign n13291 = n13259[63:62]; // extract
  /* TG68K_FPU_Transcendental.vhd:1425:49  */
  assign n13292 = n13237 ? n13291 : n13287;
  /* TG68K_FPU_Transcendental.vhd:1423:41  */
  assign n13294 = trans_state == 3'b110;
  /* TG68K_FPU_Transcendental.vhd:1460:71  */
  assign n13295 = {result_sign, result_exp};
  /* TG68K_FPU_Transcendental.vhd:1460:84  */
  assign n13296 = {n13295, result_mant};
  /* TG68K_FPU_Transcendental.vhd:1458:41  */
  assign n13298 = trans_state == 3'b111;
  assign n13299 = {n13298, n13294, n13232, n13097, n13095, n11257, n11167, n11124};
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13301 = n13296;
      8'b01000000: n13301 = n13636;
      8'b00100000: n13301 = n13636;
      8'b00010000: n13301 = n13636;
      8'b00001000: n13301 = n13636;
      8'b00000100: n13301 = n13636;
      8'b00000010: n13301 = n13636;
      8'b00000001: n13301 = n13636;
      default: n13301 = 80'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13305 = 1'b1;
      8'b01000000: n13305 = n13638;
      8'b00100000: n13305 = n13638;
      8'b00010000: n13305 = n13638;
      8'b00001000: n13305 = n13638;
      8'b00000100: n13305 = n13638;
      8'b00000010: n13305 = n13638;
      8'b00000001: n13305 = 1'b0;
      default: n13305 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13308 = 1'b0;
      8'b01000000: n13308 = n13640;
      8'b00100000: n13308 = n13640;
      8'b00010000: n13308 = n13640;
      8'b00001000: n13308 = n13640;
      8'b00000100: n13308 = n13640;
      8'b00000010: n13308 = n13640;
      8'b00000001: n13308 = n11115;
      default: n13308 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13312 = 1'b1;
      8'b01000000: n13312 = n13642;
      8'b00100000: n13312 = n13642;
      8'b00010000: n13312 = n13642;
      8'b00001000: n13312 = n13642;
      8'b00000100: n13312 = n13642;
      8'b00000010: n13312 = n13642;
      8'b00000001: n13312 = 1'b0;
      default: n13312 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13317 = 3'b000;
      8'b01000000: n13317 = 3'b111;
      8'b00100000: n13317 = n13219;
      8'b00010000: n13317 = 3'b110;
      8'b00001000: n13317 = n13065;
      8'b00000100: n13317 = n11249;
      8'b00000010: n13317 = n11160;
      8'b00000001: n13317 = n11118;
      default: n13317 = 3'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13319 = cordic_x;
      8'b01000000: n13319 = cordic_x;
      8'b00100000: n13319 = n13220;
      8'b00010000: n13319 = cordic_x;
      8'b00001000: n13319 = cordic_x;
      8'b00000100: n13319 = cordic_x;
      8'b00000010: n13319 = cordic_x;
      8'b00000001: n13319 = cordic_x;
      default: n13319 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13321 = cordic_y;
      8'b01000000: n13321 = cordic_y;
      8'b00100000: n13321 = n13221;
      8'b00010000: n13321 = cordic_y;
      8'b00001000: n13321 = cordic_y;
      8'b00000100: n13321 = cordic_y;
      8'b00000010: n13321 = cordic_y;
      8'b00000001: n13321 = cordic_y;
      default: n13321 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13323 = cordic_z;
      8'b01000000: n13323 = cordic_z;
      8'b00100000: n13323 = n13222;
      8'b00010000: n13323 = cordic_z;
      8'b00001000: n13323 = cordic_z;
      8'b00000100: n13323 = cordic_z;
      8'b00000010: n13323 = cordic_z;
      8'b00000001: n13323 = cordic_z;
      default: n13323 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13325 = cordic_iteration;
      8'b01000000: n13325 = cordic_iteration;
      8'b00100000: n13325 = n13223;
      8'b00010000: n13325 = cordic_iteration;
      8'b00001000: n13325 = n13066;
      8'b00000100: n13325 = cordic_iteration;
      8'b00000010: n13325 = cordic_iteration;
      8'b00000001: n13325 = cordic_iteration;
      default: n13325 = 5'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13327 = cordic_mode;
      8'b01000000: n13327 = cordic_mode;
      8'b00100000: n13327 = n13224;
      8'b00010000: n13327 = cordic_mode;
      8'b00001000: n13327 = cordic_mode;
      8'b00000100: n13327 = cordic_mode;
      8'b00000010: n13327 = cordic_mode;
      8'b00000001: n13327 = cordic_mode;
      default: n13327 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13329 = result_sign;
      8'b01000000: n13329 = result_sign;
      8'b00100000: n13329 = n13225;
      8'b00010000: n13329 = result_sign;
      8'b00001000: n13329 = n13068;
      8'b00000100: n13329 = n11250;
      8'b00000010: n13329 = n11161;
      8'b00000001: n13329 = result_sign;
      default: n13329 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13331 = result_exp;
      8'b01000000: n13331 = n13258;
      8'b00100000: n13331 = n13226;
      8'b00010000: n13331 = result_exp;
      8'b00001000: n13331 = n13070;
      8'b00000100: n13331 = n11251;
      8'b00000010: n13331 = n11163;
      8'b00000001: n13331 = result_exp;
      default: n13331 = 15'bX;
    endcase
  assign n13332 = n11164[61:0]; // extract
  assign n13333 = n11252[61:0]; // extract
  assign n13334 = n13072[61:0]; // extract
  assign n13335 = n13227[61:0]; // extract
  assign n13336 = result_mant[61:0]; // extract
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13338 = n13336;
      8'b01000000: n13338 = n13290;
      8'b00100000: n13338 = n13335;
      8'b00010000: n13338 = n13336;
      8'b00001000: n13338 = n13334;
      8'b00000100: n13338 = n13333;
      8'b00000010: n13338 = n13332;
      8'b00000001: n13338 = n13336;
      default: n13338 = 62'bX;
    endcase
  assign n13339 = n11164[63:62]; // extract
  assign n13340 = n11252[63:62]; // extract
  assign n13341 = n13072[63:62]; // extract
  assign n13342 = n13227[63:62]; // extract
  assign n13343 = result_mant[63:62]; // extract
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13345 = n13343;
      8'b01000000: n13345 = n13292;
      8'b00100000: n13345 = n13342;
      8'b00010000: n13345 = n13343;
      8'b00001000: n13345 = n13341;
      8'b00000100: n13345 = n13340;
      8'b00000010: n13345 = n13339;
      8'b00000001: n13345 = n13343;
      default: n13345 = 2'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13349 = series_term;
      8'b01000000: n13349 = series_term;
      8'b00100000: n13349 = series_term;
      8'b00010000: n13349 = series_term;
      8'b00001000: n13349 = n13073;
      8'b00000100: n13349 = series_term;
      8'b00000010: n13349 = series_term;
      8'b00000001: n13349 = series_term;
      default: n13349 = 80'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13351 = series_sum;
      8'b01000000: n13351 = series_sum;
      8'b00100000: n13351 = series_sum;
      8'b00010000: n13351 = series_sum;
      8'b00001000: n13351 = n13074;
      8'b00000100: n13351 = series_sum;
      8'b00000010: n13351 = series_sum;
      8'b00000001: n13351 = series_sum;
      default: n13351 = 80'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13353 = iteration_count;
      8'b01000000: n13353 = iteration_count;
      8'b00100000: n13353 = iteration_count;
      8'b00010000: n13353 = iteration_count;
      8'b00001000: n13353 = n13075;
      8'b00000100: n13353 = iteration_count;
      8'b00000010: n13353 = iteration_count;
      8'b00000001: n13353 = n11122;
      default: n13353 = 4'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13356 = trans_overflow;
      8'b01000000: n13356 = trans_overflow;
      8'b00100000: n13356 = trans_overflow;
      8'b00010000: n13356 = trans_overflow;
      8'b00001000: n13356 = n13076;
      8'b00000100: n13356 = trans_overflow;
      8'b00000010: n13356 = trans_overflow;
      8'b00000001: n13356 = 1'b0;
      default: n13356 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13359 = trans_underflow;
      8'b01000000: n13359 = trans_underflow;
      8'b00100000: n13359 = trans_underflow;
      8'b00010000: n13359 = trans_underflow;
      8'b00001000: n13359 = n13077;
      8'b00000100: n13359 = trans_underflow;
      8'b00000010: n13359 = trans_underflow;
      8'b00000001: n13359 = 1'b0;
      default: n13359 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13362 = trans_inexact;
      8'b01000000: n13362 = trans_inexact;
      8'b00100000: n13362 = trans_inexact;
      8'b00010000: n13362 = trans_inexact;
      8'b00001000: n13362 = n13080;
      8'b00000100: n13362 = trans_inexact;
      8'b00000010: n13362 = trans_inexact;
      8'b00000001: n13362 = 1'b0;
      default: n13362 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13365 = trans_invalid;
      8'b01000000: n13365 = trans_invalid;
      8'b00100000: n13365 = trans_invalid;
      8'b00010000: n13365 = trans_invalid;
      8'b00001000: n13365 = n13082;
      8'b00000100: n13365 = n11253;
      8'b00000010: n13365 = n11165;
      8'b00000001: n13365 = 1'b0;
      default: n13365 = 1'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13369 = exp_argument;
      8'b01000000: n13369 = exp_argument;
      8'b00100000: n13369 = exp_argument;
      8'b00010000: n13369 = exp_argument;
      8'b00001000: n13369 = n13083;
      8'b00000100: n13369 = exp_argument;
      8'b00000010: n13369 = exp_argument;
      8'b00000001: n13369 = exp_argument;
      default: n13369 = 80'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13371 = log_argument;
      8'b01000000: n13371 = log_argument;
      8'b00100000: n13371 = log_argument;
      8'b00010000: n13371 = log_argument;
      8'b00001000: n13371 = n13084;
      8'b00000100: n13371 = n11255;
      8'b00000010: n13371 = log_argument;
      8'b00000001: n13371 = log_argument;
      default: n13371 = 80'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13373 = x_squared;
      8'b01000000: n13373 = x_squared;
      8'b00100000: n13373 = x_squared;
      8'b00010000: n13373 = x_squared;
      8'b00001000: n13373 = n13085;
      8'b00000100: n13373 = x_squared;
      8'b00000010: n13373 = x_squared;
      8'b00000001: n13373 = x_squared;
      default: n13373 = 128'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13375 = x_cubed;
      8'b01000000: n13375 = x_cubed;
      8'b00100000: n13375 = x_cubed;
      8'b00010000: n13375 = x_cubed;
      8'b00001000: n13375 = n13086;
      8'b00000100: n13375 = x_cubed;
      8'b00000010: n13375 = x_cubed;
      8'b00000001: n13375 = x_cubed;
      default: n13375 = 128'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13377 = x_fifth;
      8'b01000000: n13377 = x_fifth;
      8'b00100000: n13377 = x_fifth;
      8'b00010000: n13377 = x_fifth;
      8'b00001000: n13377 = n13087;
      8'b00000100: n13377 = x_fifth;
      8'b00000010: n13377 = x_fifth;
      8'b00000001: n13377 = x_fifth;
      default: n13377 = 128'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13379 = x3_div6;
      8'b01000000: n13379 = x3_div6;
      8'b00100000: n13379 = x3_div6;
      8'b00010000: n13379 = x3_div6;
      8'b00001000: n13379 = n13088;
      8'b00000100: n13379 = x3_div6;
      8'b00000010: n13379 = x3_div6;
      8'b00000001: n13379 = x3_div6;
      default: n13379 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13381 = cordic_shift_x;
      8'b01000000: n13381 = cordic_shift_x;
      8'b00100000: n13381 = n13228;
      8'b00010000: n13381 = cordic_shift_x;
      8'b00001000: n13381 = cordic_shift_x;
      8'b00000100: n13381 = cordic_shift_x;
      8'b00000010: n13381 = cordic_shift_x;
      8'b00000001: n13381 = cordic_shift_x;
      default: n13381 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13383 = cordic_shift_y;
      8'b01000000: n13383 = cordic_shift_y;
      8'b00100000: n13383 = n13229;
      8'b00010000: n13383 = cordic_shift_y;
      8'b00001000: n13383 = cordic_shift_y;
      8'b00000100: n13383 = cordic_shift_y;
      8'b00000010: n13383 = cordic_shift_y;
      8'b00000001: n13383 = cordic_shift_y;
      default: n13383 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13385 = cordic_atan_val;
      8'b01000000: n13385 = cordic_atan_val;
      8'b00100000: n13385 = n13230;
      8'b00010000: n13385 = cordic_atan_val;
      8'b00001000: n13385 = cordic_atan_val;
      8'b00000100: n13385 = cordic_atan_val;
      8'b00000010: n13385 = cordic_atan_val;
      8'b00000001: n13385 = cordic_atan_val;
      default: n13385 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13387 = x5_div120;
      8'b01000000: n13387 = x5_div120;
      8'b00100000: n13387 = x5_div120;
      8'b00010000: n13387 = x5_div120;
      8'b00001000: n13387 = n13089;
      8'b00000100: n13387 = x5_div120;
      8'b00000010: n13387 = x5_div120;
      8'b00000001: n13387 = x5_div120;
      default: n13387 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13389 = x_n;
      8'b01000000: n13389 = x_n;
      8'b00100000: n13389 = x_n;
      8'b00010000: n13389 = x_n;
      8'b00001000: n13389 = n13090;
      8'b00000100: n13389 = x_n;
      8'b00000010: n13389 = x_n;
      8'b00000001: n13389 = x_n;
      default: n13389 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13391 = a_div_x_n;
      8'b01000000: n13391 = a_div_x_n;
      8'b00100000: n13391 = a_div_x_n;
      8'b00010000: n13391 = a_div_x_n;
      8'b00001000: n13391 = n13091;
      8'b00000100: n13391 = a_div_x_n;
      8'b00000010: n13391 = a_div_x_n;
      8'b00000001: n13391 = a_div_x_n;
      default: n13391 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13393 = x_next;
      8'b01000000: n13393 = x_next;
      8'b00100000: n13393 = x_next;
      8'b00010000: n13393 = x_next;
      8'b00001000: n13393 = n13092;
      8'b00000100: n13393 = x_next;
      8'b00000010: n13393 = x_next;
      8'b00000001: n13393 = x_next;
      default: n13393 = 64'bX;
    endcase
  /* TG68K_FPU_Transcendental.vhd:232:33  */
  always @*
    case (n13299)
      8'b10000000: n13395 = final_mant;
      8'b01000000: n13395 = final_mant;
      8'b00100000: n13395 = final_mant;
      8'b00010000: n13395 = final_mant;
      8'b00001000: n13395 = n13093;
      8'b00000100: n13395 = final_mant;
      8'b00000010: n13395 = final_mant;
      8'b00000001: n13395 = final_mant;
      default: n13395 = 64'bX;
    endcase
  assign n13408 = {n13345, n13338};
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13515 = clkena ? n13317 : trans_state;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13516 <= 3'b000;
    else
      n13516 <= n13515;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13517 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13518 = clkena & n13517;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13519 = n13518 ? n13319 : cordic_x;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13520 <= n13519;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13521 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13522 = clkena & n13521;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13523 = n13522 ? n13321 : cordic_y;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13524 <= n13523;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13525 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13526 = clkena & n13525;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13527 = n13526 ? n13323 : cordic_z;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13528 <= n13527;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13529 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13530 = clkena & n13529;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13531 = n13530 ? n13325 : cordic_iteration;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13532 <= n13531;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13533 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13534 = clkena & n13533;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13535 = n13534 ? n13327 : cordic_mode;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13536 <= n13535;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13537 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13538 = clkena & n13537;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13539 = n13538 ? n13329 : result_sign;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13540 <= n13539;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13541 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13542 = clkena & n13541;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13543 = n13542 ? n13331 : result_exp;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13544 <= n13543;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13545 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13546 = clkena & n13545;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13547 = n13546 ? n13408 : result_mant;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13548 <= n13547;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13553 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13554 = clkena & n13553;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13555 = n13554 ? n13349 : series_term;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13556 <= n13555;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13557 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13558 = clkena & n13557;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13559 = n13558 ? n13351 : series_sum;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13560 <= n13559;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13561 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13562 = clkena & n13561;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13563 = n13562 ? n13353 : iteration_count;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13564 <= n13563;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13565 = clkena ? n13356 : trans_overflow;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13566 <= 1'b0;
    else
      n13566 <= n13565;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13567 = clkena ? n13359 : trans_underflow;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13568 <= 1'b0;
    else
      n13568 <= n13567;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13569 = clkena ? n13362 : trans_inexact;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13570 <= 1'b0;
    else
      n13570 <= n13569;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13571 = clkena ? n13365 : trans_invalid;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13572 <= 1'b0;
    else
      n13572 <= n13571;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13577 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13578 = clkena & n13577;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13579 = n13578 ? n13369 : exp_argument;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13580 <= n13579;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13581 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13582 = clkena & n13581;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13583 = n13582 ? n13371 : log_argument;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13584 <= n13583;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13586 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13587 = clkena & n13586;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13588 = n13587 ? n13373 : x_squared;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13589 <= n13588;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13590 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13591 = clkena & n13590;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13592 = n13591 ? n13375 : x_cubed;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13593 <= n13592;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13594 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13595 = clkena & n13594;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13596 = n13595 ? n13377 : x_fifth;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13597 <= n13596;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13598 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13599 = clkena & n13598;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13600 = n13599 ? n13379 : x3_div6;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13601 <= n13600;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13602 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13603 = clkena & n13602;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13604 = n13603 ? n13381 : cordic_shift_x;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13605 <= n13604;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13606 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13607 = clkena & n13606;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13608 = n13607 ? n13383 : cordic_shift_y;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13609 <= n13608;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13610 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13611 = clkena & n13610;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13612 = n13611 ? n13385 : cordic_atan_val;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13613 <= n13612;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13614 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13615 = clkena & n13614;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13616 = n13615 ? n13387 : x5_div120;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13617 <= n13616;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13619 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13620 = clkena & n13619;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13621 = n13620 ? n13389 : x_n;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13622 <= n13621;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13623 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13624 = clkena & n13623;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13625 = n13624 ? n13391 : a_div_x_n;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13626 <= n13625;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13627 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13628 = clkena & n13627;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13629 = n13628 ? n13393 : x_next;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13630 <= n13629;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13631 = ~n11111;
  /* TG68K_FPU_Transcendental.vhd:217:9  */
  assign n13632 = clkena & n13631;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13633 = n13632 ? n13395 : final_mant;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk)
    n13634 <= n13633;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13635 = clkena ? n13301 : n13636;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13636 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n13636 <= n13635;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13637 = clkena ? n13305 : n13638;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13638 <= 1'b0;
    else
      n13638 <= n13637;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13639 = clkena ? n13308 : n13640;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13640 <= 1'b0;
    else
      n13640 <= n13639;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  assign n13641 = clkena ? n13312 : n13642;
  /* TG68K_FPU_Transcendental.vhd:230:17  */
  always @(posedge clk or posedge n11111)
    if (n11111)
      n13642 <= 1'b0;
    else
      n13642 <= n13641;
  /* TG68K_FPU_Transcendental.vhd:1369:118  */
  reg [63:0] n13643[15:0] ; // memory
  initial begin
    n13643[15] = 64'b0000000000000001111111111111111111111111111111111111111111111111;
    n13643[14] = 64'b0000000000000011111111111111111111111111111111111111111010101011;
    n13643[13] = 64'b0000000000000111111111111111111111111111111111111111010101010101;
    n13643[12] = 64'b0000000000001111111111111111111111111111111110101010101010101011;
    n13643[11] = 64'b0000000000011111111111111111111111111110101010101010101010101011;
    n13643[10] = 64'b0000000000111111111111111111111111110101010101011010101010101011;
    n13643[9] = 64'b0000000001111111111111111111110101010101010110101011101110011101;
    n13643[8] = 64'b0000000011111111111111111010101010101011010101010101011101101011;
    n13643[7] = 64'b0000000111111111111111010101010101011011101110111001011101110110;
    n13643[6] = 64'b0000001111111111111010101010101101110111010101110011101010111010;
    n13643[5] = 64'b0000011111111111010101010110111011101010010111110111101001011110;
    n13643[4] = 64'b0000111111111010101011011110100011010101101110001111000010111011;
    n13643[3] = 64'b0001111111010101101110101001101010101100001011110110101011000101;
    n13643[2] = 64'b0011111010110110111010111111001011011001001001111101101011010100;
    n13643[1] = 64'b0111011010110001100111000001010110000110010100001001111100100110;
    n13643[0] = 64'b1100100100001111110110101010001000100001011010001100001000110101;
    end
  assign n13645 = n13643[n13151];
  /* TG68K_FPU_Transcendental.vhd:1369:118  */
endmodule

module tg68k_fpu_alu
  (input  clk,
   input  nreset,
   input  clkena,
   input  start_operation,
   input  [6:0] operation_code,
   input  [1:0] rounding_mode,
   input  [79:0] operand_a,
   input  [79:0] operand_b,
   output [79:0] result,
   output result_valid,
   output overflow,
   output underflow,
   output inexact,
   output invalid,
   output divide_by_zero,
   output [7:0] quotient_byte,
   output operation_busy,
   output operation_done);
  wire sign_a;
  wire sign_b;
  wire sign_result;
  wire [14:0] exp_a;
  wire [14:0] exp_b;
  wire [14:0] exp_result;
  wire [63:0] mant_a;
  wire [63:0] mant_b;
  wire [63:0] mant_result;
  reg [2:0] alu_state;
  wire [64:0] mant_sum;
  wire [64:0] mant_a_aligned;
  wire [64:0] mant_b_aligned;
  wire [14:0] exp_larger;
  wire guard_bit;
  wire round_bit;
  wire sticky_bit;
  wire [127:0] mult_result;
  reg [7:0] fmod_quotient;
  wire is_zero_a;
  wire is_zero_b;
  wire is_inf_a;
  wire is_inf_b;
  wire is_nan_a;
  wire is_nan_b;
  wire is_denorm_a;
  wire is_denorm_b;
  wire is_snan_a;
  wire is_snan_b;
  wire flags_overflow;
  wire flags_underflow;
  wire flags_inexact;
  wire flags_invalid;
  wire flags_div_by_zero;
  wire [14:0] n7356;
  wire n7358;
  wire [63:0] n7359;
  wire n7361;
  wire n7364;
  wire n7367;
  wire [14:0] n7368;
  wire n7370;
  wire [63:0] n7371;
  wire n7373;
  wire n7374;
  wire n7375;
  wire [61:0] n7376;
  wire n7378;
  wire n7379;
  wire n7382;
  wire n7388;
  wire n7391;
  wire n7393;
  wire n7397;
  wire n7399;
  wire n7401;
  wire n7405;
  wire n7407;
  wire n7409;
  wire n7411;
  wire n7413;
  wire [14:0] n7416;
  wire n7418;
  wire [63:0] n7419;
  wire n7421;
  wire n7424;
  wire n7427;
  wire [14:0] n7428;
  wire n7430;
  wire [63:0] n7431;
  wire n7433;
  wire n7434;
  wire n7435;
  wire [61:0] n7436;
  wire n7438;
  wire n7439;
  wire n7442;
  wire n7448;
  wire n7451;
  wire n7453;
  wire n7457;
  wire n7459;
  wire n7461;
  wire n7465;
  wire n7467;
  wire n7469;
  wire n7471;
  wire n7473;
  wire n7481;
  wire n7485;
  wire [2:0] n7488;
  wire n7490;
  wire n7492;
  wire n7493;
  wire [14:0] n7494;
  wire [63:0] n7495;
  wire n7496;
  wire [14:0] n7497;
  wire [63:0] n7498;
  wire n7500;
  wire n7501;
  wire [14:0] n7502;
  wire [63:0] n7503;
  wire n7505;
  wire n7506;
  wire n7507;
  wire n7508;
  wire n7509;
  wire [14:0] n7510;
  wire [63:0] n7511;
  wire n7513;
  wire n7514;
  wire n7515;
  wire n7516;
  wire n7517;
  wire n7518;
  wire n7519;
  wire [14:0] n7521;
  wire [63:0] n7523;
  wire [2:0] n7526;
  wire n7527;
  wire [14:0] n7528;
  wire [63:0] n7529;
  wire [2:0] n7531;
  wire n7532;
  wire [14:0] n7533;
  wire [63:0] n7534;
  wire [2:0] n7536;
  wire n7538;
  wire n7540;
  wire n7542;
  wire n7543;
  wire n7545;
  wire n7546;
  wire n7547;
  wire [30:0] n7548;
  wire [31:0] n7549;
  wire [31:0] n7551;
  wire [31:0] n7553;
  wire [31:0] n7555;
  wire [30:0] n7556;
  wire [14:0] n7557;
  wire [1:0] n7558;
  wire n7560;
  wire [1:0] n7561;
  wire n7563;
  wire [1:0] n7564;
  wire n7566;
  wire [63:0] n7569;
  wire [63:0] n7571;
  wire [63:0] n7573;
  wire n7574;
  wire [62:0] n7575;
  wire [63:0] n7576;
  wire [63:0] n7577;
  wire [63:0] n7578;
  wire [14:0] n7580;
  wire [63:0] n7582;
  wire n7584;
  wire [14:0] n7587;
  wire [63:0] n7589;
  wire n7590;
  wire [14:0] n7593;
  wire [63:0] n7595;
  wire n7596;
  wire n7598;
  wire n7601;
  wire n7602;
  wire n7603;
  wire n7605;
  wire n7606;
  wire n7607;
  wire n7609;
  wire [63:0] n7612;
  wire n7614;
  wire n7615;
  wire n7616;
  wire n7617;
  wire n7618;
  wire n7619;
  wire n7621;
  wire [64:0] n7623;
  wire [64:0] n7625;
  wire [64:0] n7626;
  wire n7628;
  wire [64:0] n7630;
  wire [64:0] n7632;
  wire [64:0] n7633;
  wire n7634;
  wire [64:0] n7635;
  wire n7636;
  wire [64:0] n7637;
  wire [64:0] n7638;
  wire n7639;
  wire [64:0] n7640;
  wire n7641;
  wire [64:0] n7642;
  wire n7643;
  wire [64:0] n7646;
  wire [14:0] n7647;
  wire n7649;
  wire [64:0] n7654;
  wire [14:0] n7655;
  wire [30:0] n7656;
  wire [64:0] n7657;
  wire [64:0] n7660;
  wire [64:0] n7663;
  wire [14:0] n7664;
  wire n7666;
  wire [64:0] n7671;
  wire [14:0] n7672;
  wire [30:0] n7673;
  wire [64:0] n7674;
  wire [64:0] n7677;
  wire [64:0] n7680;
  wire [64:0] n7681;
  wire [14:0] n7682;
  wire n7684;
  wire [64:0] n7685;
  wire n7686;
  wire [64:0] n7687;
  wire [64:0] n7688;
  wire n7689;
  wire [64:0] n7690;
  wire n7691;
  wire [64:0] n7692;
  wire n7693;
  wire [14:0] n7695;
  wire [63:0] n7696;
  wire n7697;
  wire n7698;
  wire [14:0] n7700;
  wire [62:0] n7701;
  wire [63:0] n7703;
  wire [63:0] n7704;
  wire [14:0] n7705;
  wire [63:0] n7706;
  wire [14:0] n7707;
  wire [63:0] n7708;
  wire n7709;
  wire [14:0] n7710;
  wire [63:0] n7711;
  wire [64:0] n7712;
  wire [64:0] n7715;
  wire [64:0] n7716;
  wire [14:0] n7718;
  wire n7720;
  wire [14:0] n7721;
  wire [63:0] n7722;
  wire [64:0] n7723;
  wire [64:0] n7726;
  wire [64:0] n7727;
  wire [14:0] n7728;
  wire n7730;
  wire [14:0] n7731;
  wire [63:0] n7732;
  wire [64:0] n7733;
  wire [64:0] n7736;
  wire [64:0] n7737;
  wire [14:0] n7738;
  wire n7740;
  wire [14:0] n7742;
  wire [63:0] n7744;
  wire [64:0] n7745;
  wire [64:0] n7748;
  wire [64:0] n7749;
  wire [14:0] n7750;
  wire n7752;
  wire [14:0] n7754;
  wire [63:0] n7756;
  wire [64:0] n7757;
  wire [64:0] n7760;
  wire [64:0] n7761;
  wire [14:0] n7762;
  wire n7764;
  wire [14:0] n7766;
  wire [63:0] n7767;
  wire [64:0] n7768;
  wire [64:0] n7771;
  wire [64:0] n7772;
  wire [14:0] n7773;
  wire n7775;
  wire n7777;
  wire [14:0] n7779;
  wire [63:0] n7781;
  wire [64:0] n7782;
  wire [64:0] n7785;
  wire [64:0] n7786;
  wire [14:0] n7787;
  wire n7789;
  wire n7791;
  wire n7792;
  wire n7793;
  wire n7794;
  wire n7796;
  wire [63:0] n7799;
  wire n7801;
  wire n7802;
  wire n7803;
  wire n7804;
  wire n7805;
  wire n7806;
  wire n7807;
  wire n7808;
  wire n7810;
  wire [64:0] n7812;
  wire [64:0] n7814;
  wire [64:0] n7815;
  wire n7817;
  wire [64:0] n7819;
  wire [64:0] n7821;
  wire [64:0] n7822;
  wire n7823;
  wire n7824;
  wire [64:0] n7825;
  wire [64:0] n7826;
  wire n7827;
  wire n7828;
  wire [64:0] n7829;
  wire [64:0] n7830;
  wire n7831;
  wire [64:0] n7832;
  wire n7833;
  wire [64:0] n7836;
  wire [14:0] n7837;
  wire n7839;
  wire [64:0] n7841;
  wire [14:0] n7842;
  wire [30:0] n7843;
  wire [64:0] n7844;
  wire [64:0] n7846;
  wire [64:0] n7849;
  wire [14:0] n7850;
  wire n7852;
  wire [64:0] n7854;
  wire [14:0] n7855;
  wire [30:0] n7856;
  wire [64:0] n7857;
  wire [64:0] n7859;
  wire [64:0] n7861;
  wire [64:0] n7862;
  wire [14:0] n7863;
  wire n7864;
  wire [64:0] n7865;
  wire n7866;
  wire [64:0] n7867;
  wire [64:0] n7868;
  wire n7869;
  wire n7870;
  wire [64:0] n7871;
  wire n7872;
  wire [64:0] n7873;
  wire n7874;
  wire [14:0] n7876;
  wire [63:0] n7877;
  wire n7878;
  wire n7879;
  wire [14:0] n7881;
  wire [62:0] n7882;
  wire [63:0] n7884;
  wire [63:0] n7885;
  wire [14:0] n7886;
  wire [63:0] n7887;
  wire [14:0] n7888;
  wire [63:0] n7889;
  wire n7890;
  wire [14:0] n7891;
  wire [63:0] n7892;
  wire [64:0] n7893;
  wire [64:0] n7895;
  wire [64:0] n7896;
  wire [14:0] n7898;
  wire n7899;
  wire [14:0] n7900;
  wire [63:0] n7901;
  wire [64:0] n7902;
  wire [64:0] n7904;
  wire [64:0] n7905;
  wire [14:0] n7906;
  wire n7907;
  wire [14:0] n7908;
  wire [63:0] n7909;
  wire [64:0] n7910;
  wire [64:0] n7912;
  wire [64:0] n7913;
  wire [14:0] n7914;
  wire n7915;
  wire [14:0] n7917;
  wire [63:0] n7919;
  wire [64:0] n7920;
  wire [64:0] n7922;
  wire [64:0] n7923;
  wire [14:0] n7924;
  wire n7925;
  wire [14:0] n7927;
  wire [63:0] n7929;
  wire [64:0] n7930;
  wire [64:0] n7932;
  wire [64:0] n7933;
  wire [14:0] n7934;
  wire n7935;
  wire [14:0] n7937;
  wire [63:0] n7938;
  wire [64:0] n7939;
  wire [64:0] n7941;
  wire [64:0] n7942;
  wire [14:0] n7943;
  wire n7944;
  wire n7946;
  wire [14:0] n7948;
  wire [63:0] n7950;
  wire [64:0] n7951;
  wire [64:0] n7953;
  wire [64:0] n7954;
  wire [14:0] n7955;
  wire n7957;
  wire n7959;
  wire n7960;
  wire n7961;
  wire n7962;
  wire n7963;
  wire n7964;
  wire n7965;
  wire n7966;
  wire [14:0] n7967;
  wire [14:0] n7969;
  wire [127:0] n7970;
  wire [127:0] n7971;
  wire [127:0] n7972;
  wire n7973;
  wire [14:0] n7975;
  wire [63:0] n7976;
  wire [63:0] n7977;
  wire [14:0] n7978;
  wire [63:0] n7979;
  wire [61:0] n7980;
  wire n7982;
  wire n7984;
  wire [14:0] n7986;
  wire [63:0] n7988;
  wire [127:0] n7989;
  wire n7990;
  wire [14:0] n7992;
  wire [63:0] n7994;
  wire [127:0] n7995;
  wire n7996;
  wire n7998;
  wire [14:0] n8000;
  wire [63:0] n8002;
  wire [127:0] n8003;
  wire n8004;
  wire n8006;
  wire n8008;
  wire [14:0] n8010;
  wire [63:0] n8012;
  wire [127:0] n8013;
  wire n8014;
  wire n8016;
  wire n8018;
  wire n8019;
  wire n8020;
  wire n8021;
  wire n8022;
  wire n8023;
  wire n8024;
  wire n8025;
  wire n8026;
  wire n8027;
  wire n8028;
  wire n8033;
  wire [31:0] n8034;
  wire n8036;
  wire [14:0] n8038;
  wire [14:0] n8040;
  wire n8041;
  wire n8042;
  wire [14:0] n8044;
  wire [63:0] n8046;
  wire n8050;
  wire [14:0] n8051;
  wire [14:0] n8053;
  wire [31:0] n8054;
  wire n8056;
  wire [63:0] n8058;
  wire [31:0] n8059;
  wire [63:0] n8060;
  wire [63:0] n8061;
  wire [47:0] n8062;
  wire n8064;
  wire [63:0] n8066;
  wire [47:0] n8067;
  wire [63:0] n8068;
  wire [63:0] n8069;
  wire [62:0] n8070;
  wire [63:0] n8071;
  wire [63:0] n8072;
  wire [63:0] n8073;
  wire [63:0] n8074;
  wire [14:0] n8076;
  wire [63:0] n8078;
  wire n8080;
  wire [14:0] n8082;
  wire [63:0] n8084;
  wire n8085;
  wire [14:0] n8087;
  wire [63:0] n8089;
  wire n8090;
  wire n8091;
  wire [14:0] n8092;
  wire [63:0] n8093;
  wire n8095;
  wire n8096;
  wire n8097;
  wire [14:0] n8099;
  wire [63:0] n8101;
  wire n8103;
  wire n8104;
  wire n8106;
  wire n8108;
  wire [14:0] n8110;
  wire [63:0] n8112;
  wire n8114;
  wire n8115;
  wire n8117;
  wire n8118;
  wire n8120;
  wire [14:0] n8122;
  wire [63:0] n8124;
  wire n8126;
  wire n8127;
  wire n8129;
  wire n8130;
  wire n8132;
  wire n8134;
  wire n8135;
  wire n8136;
  wire n8138;
  wire n8139;
  wire n8140;
  wire n8142;
  wire n8145;
  wire n8146;
  wire n8147;
  wire n8150;
  wire n8151;
  wire n8152;
  wire n8155;
  wire n8156;
  wire n8157;
  wire n8158;
  wire [78:0] n8159;
  wire [78:0] n8160;
  wire n8161;
  wire n8162;
  wire n8165;
  wire n8167;
  wire n8168;
  wire n8169;
  wire n8171;
  wire n8173;
  wire n8176;
  wire n8178;
  wire n8180;
  wire n8181;
  wire n8183;
  wire n8185;
  wire n8186;
  wire n8187;
  wire [14:0] n8190;
  wire [63:0] n8193;
  wire [30:0] n8194;
  wire [31:0] n8195;
  wire [31:0] n8197;
  wire n8199;
  wire n8201;
  wire [31:0] n8203;
  wire n8205;
  wire n8207;
  wire n8208;
  wire [31:0] n8210;
  wire n8212;
  wire n8214;
  wire n8215;
  wire [31:0] n8217;
  wire n8219;
  wire n8221;
  wire n8222;
  wire [31:0] n8224;
  wire n8226;
  wire n8228;
  wire n8229;
  wire [31:0] n8231;
  wire n8233;
  wire n8235;
  wire n8236;
  wire [31:0] n8238;
  wire n8240;
  wire n8242;
  wire n8243;
  wire [31:0] n8245;
  wire n8247;
  wire n8249;
  wire n8250;
  wire [31:0] n8252;
  wire n8254;
  wire n8256;
  wire n8257;
  wire [31:0] n8259;
  wire n8261;
  wire n8263;
  wire n8264;
  wire [31:0] n8266;
  wire n8268;
  wire n8270;
  wire n8271;
  wire [31:0] n8273;
  wire n8275;
  wire n8277;
  wire n8278;
  wire [31:0] n8280;
  wire n8282;
  wire n8284;
  wire n8285;
  wire [31:0] n8287;
  wire n8289;
  wire n8291;
  wire n8292;
  wire [31:0] n8294;
  wire n8296;
  wire n8298;
  wire n8299;
  wire [31:0] n8301;
  wire n8303;
  wire n8305;
  wire n8306;
  wire [31:0] n8308;
  wire n8310;
  wire n8312;
  wire n8313;
  wire [31:0] n8315;
  wire n8317;
  wire n8319;
  wire n8320;
  wire [31:0] n8322;
  wire n8324;
  wire n8326;
  wire n8327;
  wire [31:0] n8329;
  wire n8331;
  wire n8333;
  wire n8334;
  wire [31:0] n8336;
  wire n8338;
  wire n8340;
  wire n8341;
  wire [31:0] n8343;
  wire n8345;
  wire n8347;
  wire n8348;
  wire [31:0] n8350;
  wire n8352;
  wire n8354;
  wire n8355;
  wire [31:0] n8357;
  wire n8359;
  wire n8361;
  wire n8362;
  wire [31:0] n8364;
  wire n8366;
  wire n8368;
  wire n8369;
  wire [31:0] n8371;
  wire n8373;
  wire n8375;
  wire n8376;
  wire [31:0] n8378;
  wire n8380;
  wire n8382;
  wire n8383;
  wire [31:0] n8385;
  wire n8387;
  wire n8389;
  wire n8390;
  wire [31:0] n8392;
  wire n8394;
  wire n8396;
  wire n8397;
  wire [31:0] n8399;
  wire n8401;
  wire n8403;
  wire n8404;
  wire [31:0] n8406;
  wire n8408;
  wire n8410;
  wire n8411;
  wire [31:0] n8413;
  wire n8415;
  wire n8417;
  wire n8418;
  wire [31:0] n8420;
  wire n8422;
  wire n8424;
  wire n8425;
  wire [31:0] n8427;
  wire n8429;
  wire n8431;
  wire n8432;
  wire [31:0] n8434;
  wire n8436;
  wire n8438;
  wire n8439;
  wire [31:0] n8441;
  wire n8443;
  wire n8445;
  wire n8446;
  wire [31:0] n8448;
  wire n8450;
  wire n8452;
  wire n8453;
  wire [31:0] n8455;
  wire n8457;
  wire n8459;
  wire n8460;
  wire [31:0] n8462;
  wire n8464;
  wire n8466;
  wire n8467;
  wire [31:0] n8469;
  wire n8471;
  wire n8473;
  wire n8474;
  wire [31:0] n8476;
  wire n8478;
  wire n8480;
  wire n8481;
  wire [31:0] n8483;
  wire n8485;
  wire n8487;
  wire n8488;
  wire [31:0] n8490;
  wire n8492;
  wire n8494;
  wire n8495;
  wire [31:0] n8497;
  wire n8499;
  wire n8501;
  wire n8502;
  wire [31:0] n8504;
  wire n8506;
  wire n8508;
  wire n8509;
  wire [31:0] n8511;
  wire n8513;
  wire n8515;
  wire n8516;
  wire [31:0] n8518;
  wire n8520;
  wire n8522;
  wire n8523;
  wire [31:0] n8525;
  wire n8527;
  wire n8529;
  wire n8530;
  wire [31:0] n8532;
  wire n8534;
  wire n8536;
  wire n8537;
  wire [31:0] n8539;
  wire n8541;
  wire n8543;
  wire n8544;
  wire [31:0] n8546;
  wire n8548;
  wire n8550;
  wire n8551;
  wire [31:0] n8553;
  wire n8555;
  wire n8557;
  wire n8558;
  wire [31:0] n8560;
  wire n8562;
  wire n8564;
  wire n8565;
  wire [31:0] n8567;
  wire n8569;
  wire n8571;
  wire n8572;
  wire [31:0] n8574;
  wire n8576;
  wire n8578;
  wire n8579;
  wire [31:0] n8581;
  wire n8583;
  wire n8585;
  wire n8586;
  wire [31:0] n8588;
  wire n8590;
  wire n8592;
  wire n8593;
  wire [31:0] n8595;
  wire n8597;
  wire n8599;
  wire n8600;
  wire [31:0] n8602;
  wire n8604;
  wire n8606;
  wire n8607;
  wire [31:0] n8609;
  wire n8611;
  wire n8613;
  wire n8614;
  wire [31:0] n8616;
  wire n8618;
  wire n8620;
  wire n8621;
  wire [31:0] n8623;
  wire n8625;
  wire n8627;
  wire n8628;
  wire [31:0] n8630;
  wire n8632;
  wire n8634;
  wire n8635;
  wire [31:0] n8637;
  wire n8639;
  wire n8641;
  wire n8642;
  wire n8643;
  wire [63:0] n8644;
  wire [63:0] n8645;
  wire [63:0] n8646;
  wire [14:0] n8647;
  wire [63:0] n8648;
  wire n8650;
  wire [14:0] n8653;
  wire [63:0] n8655;
  wire n8656;
  wire [14:0] n8659;
  wire [63:0] n8661;
  wire n8662;
  wire n8665;
  wire [14:0] n8667;
  wire [63:0] n8669;
  wire n8670;
  wire n8672;
  wire n8675;
  wire n8677;
  wire [30:0] n8678;
  wire [31:0] n8679;
  wire [31:0] n8681;
  wire n8683;
  wire n8685;
  wire [31:0] n8687;
  wire n8689;
  wire n8691;
  wire n8692;
  wire [31:0] n8694;
  wire n8696;
  wire n8698;
  wire n8699;
  wire [31:0] n8701;
  wire n8703;
  wire n8705;
  wire n8706;
  wire [31:0] n8708;
  wire n8710;
  wire n8712;
  wire n8713;
  wire [31:0] n8715;
  wire n8717;
  wire n8719;
  wire n8720;
  wire [31:0] n8722;
  wire n8724;
  wire n8726;
  wire n8727;
  wire [31:0] n8729;
  wire n8731;
  wire n8733;
  wire n8734;
  wire [31:0] n8736;
  wire n8738;
  wire n8740;
  wire n8741;
  wire [31:0] n8743;
  wire n8745;
  wire n8747;
  wire n8748;
  wire [31:0] n8750;
  wire n8752;
  wire n8754;
  wire n8755;
  wire [31:0] n8757;
  wire n8759;
  wire n8761;
  wire n8762;
  wire [31:0] n8764;
  wire n8766;
  wire n8768;
  wire n8769;
  wire [31:0] n8771;
  wire n8773;
  wire n8775;
  wire n8776;
  wire [31:0] n8778;
  wire n8780;
  wire n8782;
  wire n8783;
  wire [31:0] n8785;
  wire n8787;
  wire n8789;
  wire n8790;
  wire [31:0] n8792;
  wire n8794;
  wire n8796;
  wire n8797;
  wire [31:0] n8799;
  wire n8801;
  wire n8803;
  wire n8804;
  wire [31:0] n8806;
  wire n8808;
  wire n8810;
  wire n8811;
  wire [31:0] n8813;
  wire n8815;
  wire n8817;
  wire n8818;
  wire [31:0] n8820;
  wire n8822;
  wire n8824;
  wire n8825;
  wire [31:0] n8827;
  wire n8829;
  wire n8831;
  wire n8832;
  wire [31:0] n8834;
  wire n8836;
  wire n8838;
  wire n8839;
  wire [31:0] n8841;
  wire n8843;
  wire n8845;
  wire n8846;
  wire [31:0] n8848;
  wire n8850;
  wire n8852;
  wire n8853;
  wire [31:0] n8855;
  wire n8857;
  wire n8859;
  wire n8860;
  wire [31:0] n8862;
  wire n8864;
  wire n8866;
  wire n8867;
  wire [31:0] n8869;
  wire n8871;
  wire n8873;
  wire n8874;
  wire [31:0] n8876;
  wire n8878;
  wire n8880;
  wire n8881;
  wire [31:0] n8883;
  wire n8885;
  wire n8887;
  wire n8888;
  wire [31:0] n8890;
  wire n8892;
  wire n8894;
  wire n8895;
  wire [31:0] n8897;
  wire n8899;
  wire n8901;
  wire n8902;
  wire [31:0] n8904;
  wire n8906;
  wire n8908;
  wire n8909;
  wire [31:0] n8911;
  wire n8913;
  wire n8915;
  wire n8916;
  wire [31:0] n8918;
  wire n8920;
  wire n8922;
  wire n8923;
  wire [31:0] n8925;
  wire n8927;
  wire n8929;
  wire n8930;
  wire [31:0] n8932;
  wire n8934;
  wire n8936;
  wire n8937;
  wire [31:0] n8939;
  wire n8941;
  wire n8943;
  wire n8944;
  wire [31:0] n8946;
  wire n8948;
  wire n8950;
  wire n8951;
  wire [31:0] n8953;
  wire n8955;
  wire n8957;
  wire n8958;
  wire [31:0] n8960;
  wire n8962;
  wire n8964;
  wire n8965;
  wire [31:0] n8967;
  wire n8969;
  wire n8971;
  wire n8972;
  wire [31:0] n8974;
  wire n8976;
  wire n8978;
  wire n8979;
  wire [31:0] n8981;
  wire n8983;
  wire n8985;
  wire n8986;
  wire [31:0] n8988;
  wire n8990;
  wire n8992;
  wire n8993;
  wire [31:0] n8995;
  wire n8997;
  wire n8999;
  wire n9000;
  wire [31:0] n9002;
  wire n9004;
  wire n9006;
  wire n9007;
  wire [31:0] n9009;
  wire n9011;
  wire n9013;
  wire n9014;
  wire [31:0] n9016;
  wire n9018;
  wire n9020;
  wire n9021;
  wire [31:0] n9023;
  wire n9025;
  wire n9027;
  wire n9028;
  wire [31:0] n9030;
  wire n9032;
  wire n9034;
  wire n9035;
  wire [31:0] n9037;
  wire n9039;
  wire n9041;
  wire n9042;
  wire [31:0] n9044;
  wire n9046;
  wire n9048;
  wire n9049;
  wire [31:0] n9051;
  wire n9053;
  wire n9055;
  wire n9056;
  wire [31:0] n9058;
  wire n9060;
  wire n9062;
  wire n9063;
  wire [31:0] n9065;
  wire n9067;
  wire n9069;
  wire n9070;
  wire [31:0] n9072;
  wire n9074;
  wire n9076;
  wire n9077;
  wire [31:0] n9079;
  wire n9081;
  wire n9083;
  wire n9084;
  wire [31:0] n9086;
  wire n9088;
  wire n9090;
  wire n9091;
  wire [31:0] n9093;
  wire n9095;
  wire n9097;
  wire n9098;
  wire [31:0] n9100;
  wire n9102;
  wire n9104;
  wire n9105;
  wire [31:0] n9107;
  wire n9109;
  wire n9111;
  wire n9112;
  wire [31:0] n9114;
  wire n9116;
  wire n9118;
  wire n9119;
  wire [31:0] n9121;
  wire n9123;
  wire n9125;
  wire n9126;
  wire n9127;
  wire [63:0] n9128;
  wire [63:0] n9129;
  wire [63:0] n9130;
  wire [14:0] n9132;
  wire [63:0] n9134;
  wire n9136;
  wire [14:0] n9139;
  wire [63:0] n9141;
  wire n9142;
  wire [14:0] n9145;
  wire [63:0] n9147;
  wire n9148;
  wire n9151;
  wire [14:0] n9153;
  wire [63:0] n9155;
  wire n9156;
  wire n9158;
  wire n9161;
  wire n9162;
  wire n9163;
  wire n9164;
  wire n9165;
  wire n9166;
  wire n9167;
  wire n9168;
  wire [14:0] n9169;
  wire [14:0] n9171;
  wire n9172;
  wire n9173;
  wire [15:0] n9174;
  wire n9176;
  wire [31:0] n9177;
  wire [63:0] n9178;
  wire [63:0] n9180;
  wire [15:0] n9181;
  wire [63:0] n9182;
  wire [63:0] n9183;
  wire [63:0] n9185;
  wire n9187;
  wire [14:0] n9189;
  wire [15:0] n9190;
  wire n9192;
  wire [31:0] n9193;
  wire [63:0] n9194;
  wire [63:0] n9196;
  wire [15:0] n9197;
  wire [63:0] n9198;
  wire [63:0] n9199;
  wire [62:0] n9200;
  wire [63:0] n9202;
  wire [63:0] n9203;
  wire [14:0] n9204;
  wire [63:0] n9205;
  wire n9206;
  wire [14:0] n9207;
  wire [63:0] n9209;
  wire n9210;
  wire [23:0] n9212;
  wire [14:0] n9214;
  wire [63:0] n9215;
  wire [63:0] n9217;
  wire n9218;
  wire n9220;
  wire [14:0] n9222;
  wire [63:0] n9224;
  wire n9225;
  wire n9226;
  wire [14:0] n9228;
  wire [63:0] n9230;
  wire n9231;
  wire n9232;
  wire [14:0] n9234;
  wire [63:0] n9236;
  wire n9237;
  wire n9238;
  wire n9240;
  wire n9242;
  wire [14:0] n9244;
  wire [63:0] n9246;
  wire n9247;
  wire n9248;
  wire n9250;
  wire n9251;
  wire n9253;
  wire [14:0] n9255;
  wire [63:0] n9257;
  wire n9258;
  wire n9259;
  wire n9261;
  wire n9262;
  wire n9264;
  wire n9265;
  wire n9266;
  wire n9267;
  wire n9268;
  wire n9269;
  wire n9270;
  wire n9271;
  wire [14:0] n9272;
  wire [14:0] n9274;
  wire [7:0] n9275;
  wire [7:0] n9276;
  wire n9277;
  wire [63:0] n9278;
  wire [14:0] n9280;
  wire [63:0] n9282;
  wire n9284;
  wire [14:0] n9286;
  wire [63:0] n9288;
  wire n9289;
  wire n9291;
  wire [14:0] n9293;
  wire [63:0] n9295;
  wire n9296;
  wire n9298;
  wire n9300;
  wire [14:0] n9302;
  wire [63:0] n9304;
  wire n9305;
  wire n9307;
  wire n9309;
  wire n9310;
  wire n9311;
  wire n9312;
  wire n9313;
  wire [14:0] n9314;
  wire n9316;
  wire [14:0] n9317;
  wire [6:0] n9319;
  wire [7:0] n9321;
  wire [63:0] n9323;
  wire [63:0] n9324;
  wire [14:0] n9325;
  wire n9327;
  wire [63:0] n9329;
  wire [63:0] n9330;
  wire [63:0] n9331;
  wire [63:0] n9332;
  wire [7:0] n9334;
  wire [14:0] n9335;
  wire [63:0] n9336;
  wire [7:0] n9338;
  wire [14:0] n9340;
  wire [63:0] n9342;
  wire [7:0] n9343;
  wire n9345;
  wire n9347;
  wire [14:0] n9349;
  wire [63:0] n9351;
  wire [7:0] n9352;
  wire n9353;
  wire n9355;
  wire n9357;
  wire n9358;
  wire n9359;
  wire n9360;
  wire n9361;
  wire [14:0] n9362;
  wire n9364;
  wire [14:0] n9365;
  wire [6:0] n9367;
  wire [7:0] n9369;
  wire [63:0] n9371;
  wire n9372;
  wire n9373;
  wire n9374;
  wire [14:0] n9375;
  wire n9377;
  wire [63:0] n9379;
  wire n9380;
  wire n9381;
  wire n9382;
  wire [14:0] n9384;
  wire n9385;
  wire n9386;
  wire [14:0] n9387;
  wire [63:0] n9388;
  wire n9389;
  wire [14:0] n9390;
  wire [63:0] n9391;
  wire [7:0] n9393;
  wire n9394;
  wire [14:0] n9395;
  wire [63:0] n9396;
  wire [7:0] n9398;
  wire n9399;
  wire [14:0] n9401;
  wire [63:0] n9403;
  wire [7:0] n9404;
  wire n9406;
  wire n9408;
  wire [14:0] n9410;
  wire [63:0] n9412;
  wire [7:0] n9413;
  wire n9414;
  wire n9416;
  wire n9418;
  wire n9419;
  wire [30:0] n9420;
  wire [31:0] n9421;
  wire n9423;
  wire [30:0] n9424;
  wire [31:0] n9425;
  wire [31:0] n9427;
  wire [31:0] n9428;
  wire [30:0] n9429;
  wire [31:0] n9430;
  wire [31:0] n9432;
  wire [31:0] n9433;
  wire [31:0] n9434;
  wire n9437;
  wire n9439;
  wire [30:0] n9440;
  wire [14:0] n9441;
  wire [14:0] n9443;
  wire [63:0] n9445;
  wire n9447;
  wire [14:0] n9449;
  wire [63:0] n9451;
  wire n9453;
  wire n9454;
  wire [14:0] n9456;
  wire [63:0] n9458;
  wire n9459;
  wire n9460;
  wire [14:0] n9464;
  wire [63:0] n9466;
  wire n9467;
  wire n9468;
  wire n9472;
  wire [14:0] n9474;
  wire [63:0] n9476;
  wire n9477;
  wire n9478;
  wire n9480;
  wire n9484;
  wire [30:0] n9485;
  wire [31:0] n9486;
  wire [31:0] n9488;
  wire n9490;
  wire [31:0] n9492;
  wire [30:0] n9493;
  wire [14:0] n9494;
  wire [31:0] n9495;
  wire [31:0] n9497;
  wire [30:0] n9498;
  wire [14:0] n9499;
  wire n9502;
  wire [14:0] n9504;
  wire n9506;
  wire [14:0] n9508;
  wire [63:0] n9511;
  wire n9514;
  wire [14:0] n9516;
  wire [63:0] n9518;
  wire n9521;
  wire [14:0] n9523;
  wire [63:0] n9525;
  wire n9528;
  wire [14:0] n9531;
  wire [63:0] n9533;
  wire n9535;
  wire [14:0] n9537;
  wire [63:0] n9539;
  wire n9541;
  wire n9543;
  wire [14:0] n9545;
  wire [63:0] n9547;
  wire n9548;
  wire n9550;
  wire [17:0] n9551;
  reg n9555;
  reg [14:0] n9558;
  reg [63:0] n9561;
  reg [64:0] n9562;
  reg [64:0] n9565;
  reg [64:0] n9566;
  reg [14:0] n9567;
  reg [127:0] n9569;
  reg [7:0] n9570;
  reg n9571;
  reg n9572;
  reg n9573;
  reg n9575;
  reg n9576;
  wire n9580;
  wire n9582;
  wire n9584;
  wire n9585;
  wire n9587;
  wire n9588;
  wire n9589;
  wire n9590;
  wire n9592;
  wire n9598;
  wire n9600;
  wire [5:0] n9603;
  wire n9607;
  wire [5:0] n9610;
  wire n9611;
  wire [5:0] n9614;
  wire n9616;
  wire n9617;
  wire [5:0] n9619;
  wire n9623;
  wire n9625;
  wire n9626;
  wire n9628;
  wire n9629;
  wire n9630;
  wire [5:0] n9632;
  wire n9636;
  wire n9638;
  wire n9639;
  wire n9641;
  wire n9642;
  wire n9643;
  wire [5:0] n9645;
  wire n9649;
  wire n9651;
  wire n9652;
  wire n9654;
  wire n9655;
  wire n9656;
  wire [5:0] n9658;
  wire n9662;
  wire n9664;
  wire n9665;
  wire n9667;
  wire n9668;
  wire n9669;
  wire [5:0] n9671;
  wire n9675;
  wire n9677;
  wire n9678;
  wire n9680;
  wire n9681;
  wire n9682;
  wire [5:0] n9684;
  wire n9688;
  wire n9690;
  wire n9691;
  wire n9693;
  wire n9694;
  wire n9695;
  wire [5:0] n9697;
  wire n9701;
  wire n9703;
  wire n9704;
  wire n9706;
  wire n9707;
  wire n9708;
  wire [5:0] n9710;
  wire n9714;
  wire n9716;
  wire n9717;
  wire n9719;
  wire n9720;
  wire n9721;
  wire [5:0] n9723;
  wire n9727;
  wire n9729;
  wire n9730;
  wire n9732;
  wire n9733;
  wire n9734;
  wire [5:0] n9736;
  wire n9740;
  wire n9742;
  wire n9743;
  wire n9745;
  wire n9746;
  wire n9747;
  wire [5:0] n9749;
  wire n9753;
  wire n9755;
  wire n9756;
  wire n9758;
  wire n9759;
  wire n9760;
  wire [5:0] n9762;
  wire n9766;
  wire n9768;
  wire n9769;
  wire n9771;
  wire n9772;
  wire n9773;
  wire [5:0] n9775;
  wire n9779;
  wire n9781;
  wire n9782;
  wire n9784;
  wire n9785;
  wire n9786;
  wire [5:0] n9788;
  wire n9792;
  wire n9794;
  wire n9795;
  wire n9797;
  wire n9798;
  wire n9799;
  wire [5:0] n9801;
  wire n9805;
  wire n9807;
  wire n9808;
  wire n9810;
  wire n9811;
  wire n9812;
  wire [5:0] n9814;
  wire n9818;
  wire n9820;
  wire n9821;
  wire n9823;
  wire n9824;
  wire n9825;
  wire [5:0] n9827;
  wire n9831;
  wire n9833;
  wire n9834;
  wire n9836;
  wire n9837;
  wire n9838;
  wire [5:0] n9840;
  wire n9844;
  wire n9846;
  wire n9847;
  wire n9849;
  wire n9850;
  wire n9851;
  wire [5:0] n9853;
  wire n9857;
  wire n9859;
  wire n9860;
  wire n9862;
  wire n9863;
  wire n9864;
  wire [5:0] n9866;
  wire n9870;
  wire n9872;
  wire n9873;
  wire n9875;
  wire n9876;
  wire n9877;
  wire [5:0] n9879;
  wire n9883;
  wire n9885;
  wire n9886;
  wire n9888;
  wire n9889;
  wire n9890;
  wire [5:0] n9892;
  wire n9896;
  wire n9898;
  wire n9899;
  wire n9901;
  wire n9902;
  wire n9903;
  wire [5:0] n9905;
  wire n9909;
  wire n9911;
  wire n9912;
  wire n9914;
  wire n9915;
  wire n9916;
  wire [5:0] n9918;
  wire n9922;
  wire n9924;
  wire n9925;
  wire n9927;
  wire n9928;
  wire n9929;
  wire [5:0] n9931;
  wire n9935;
  wire n9937;
  wire n9938;
  wire n9940;
  wire n9941;
  wire n9942;
  wire [5:0] n9944;
  wire n9948;
  wire n9950;
  wire n9951;
  wire n9953;
  wire n9954;
  wire n9955;
  wire [5:0] n9957;
  wire n9961;
  wire n9963;
  wire n9964;
  wire n9966;
  wire n9967;
  wire n9968;
  wire [5:0] n9970;
  wire n9974;
  wire n9976;
  wire n9977;
  wire n9979;
  wire n9980;
  wire n9981;
  wire [5:0] n9983;
  wire n9987;
  wire n9989;
  wire n9990;
  wire n9992;
  wire n9993;
  wire n9994;
  wire [5:0] n9996;
  wire n10000;
  wire n10002;
  wire n10003;
  wire n10005;
  wire n10006;
  wire n10007;
  wire [5:0] n10009;
  wire n10013;
  wire n10015;
  wire n10016;
  wire n10018;
  wire n10019;
  wire n10020;
  wire [5:0] n10022;
  wire n10026;
  wire n10028;
  wire n10029;
  wire n10031;
  wire n10032;
  wire n10033;
  wire [5:0] n10035;
  wire n10039;
  wire n10041;
  wire n10042;
  wire n10044;
  wire n10045;
  wire n10046;
  wire [5:0] n10048;
  wire n10052;
  wire n10054;
  wire n10055;
  wire n10057;
  wire n10058;
  wire n10059;
  wire [5:0] n10061;
  wire n10065;
  wire n10067;
  wire n10068;
  wire n10070;
  wire n10071;
  wire n10072;
  wire [5:0] n10074;
  wire n10078;
  wire n10080;
  wire n10081;
  wire n10083;
  wire n10084;
  wire n10085;
  wire [5:0] n10087;
  wire n10091;
  wire n10093;
  wire n10094;
  wire n10096;
  wire n10097;
  wire n10098;
  wire [5:0] n10100;
  wire n10104;
  wire n10106;
  wire n10107;
  wire n10109;
  wire n10110;
  wire n10111;
  wire [5:0] n10113;
  wire n10117;
  wire n10119;
  wire n10120;
  wire n10122;
  wire n10123;
  wire n10124;
  wire [5:0] n10126;
  wire n10130;
  wire n10132;
  wire n10133;
  wire n10135;
  wire n10136;
  wire n10137;
  wire [5:0] n10139;
  wire n10143;
  wire n10145;
  wire n10146;
  wire n10148;
  wire n10149;
  wire n10150;
  wire [5:0] n10152;
  wire n10156;
  wire n10158;
  wire n10159;
  wire n10161;
  wire n10162;
  wire n10163;
  wire [5:0] n10165;
  wire n10169;
  wire n10171;
  wire n10172;
  wire n10174;
  wire n10175;
  wire n10176;
  wire [5:0] n10178;
  wire n10182;
  wire n10184;
  wire n10185;
  wire n10187;
  wire n10188;
  wire n10189;
  wire [5:0] n10191;
  wire n10195;
  wire n10197;
  wire n10198;
  wire n10200;
  wire n10201;
  wire n10202;
  wire [5:0] n10204;
  wire n10208;
  wire n10210;
  wire n10211;
  wire n10213;
  wire n10214;
  wire n10215;
  wire [5:0] n10217;
  wire n10221;
  wire n10223;
  wire n10224;
  wire n10226;
  wire n10227;
  wire n10228;
  wire [5:0] n10230;
  wire n10234;
  wire n10236;
  wire n10237;
  wire n10239;
  wire n10240;
  wire n10241;
  wire [5:0] n10243;
  wire n10247;
  wire n10249;
  wire n10250;
  wire n10252;
  wire n10253;
  wire n10254;
  wire [5:0] n10256;
  wire n10260;
  wire n10262;
  wire n10263;
  wire n10265;
  wire n10266;
  wire n10267;
  wire [5:0] n10269;
  wire n10273;
  wire n10275;
  wire n10276;
  wire n10278;
  wire n10279;
  wire n10280;
  wire [5:0] n10282;
  wire n10286;
  wire n10288;
  wire n10289;
  wire n10291;
  wire n10292;
  wire n10293;
  wire [5:0] n10295;
  wire n10299;
  wire n10301;
  wire n10302;
  wire n10304;
  wire n10305;
  wire n10306;
  wire [5:0] n10308;
  wire n10312;
  wire n10314;
  wire n10315;
  wire n10317;
  wire n10318;
  wire n10319;
  wire [5:0] n10321;
  wire n10325;
  wire n10327;
  wire n10328;
  wire n10330;
  wire n10331;
  wire n10332;
  wire [5:0] n10334;
  wire n10338;
  wire n10340;
  wire n10341;
  wire n10343;
  wire n10344;
  wire n10345;
  wire [5:0] n10347;
  wire n10351;
  wire n10353;
  wire n10354;
  wire n10356;
  wire n10357;
  wire n10358;
  wire [5:0] n10360;
  wire n10364;
  wire n10366;
  wire n10367;
  wire n10369;
  wire n10370;
  wire n10371;
  wire [5:0] n10373;
  wire n10377;
  wire n10379;
  wire n10380;
  wire n10382;
  wire n10383;
  wire n10384;
  wire [5:0] n10386;
  wire n10390;
  wire n10392;
  wire n10393;
  wire n10395;
  wire n10396;
  wire n10397;
  wire [5:0] n10399;
  wire n10403;
  wire n10405;
  wire n10406;
  wire n10408;
  wire n10409;
  wire n10410;
  wire [5:0] n10412;
  wire n10418;
  wire n10421;
  wire [31:0] n10423;
  wire n10425;
  wire n10427;
  wire n10428;
  wire n10429;
  wire n10431;
  wire n10434;
  wire n10435;
  wire n10437;
  wire n10438;
  wire n10439;
  wire n10440;
  wire n10441;
  wire n10442;
  wire n10443;
  wire n10446;
  wire n10448;
  wire n10450;
  wire n10452;
  wire n10453;
  wire n10455;
  wire n10457;
  wire n10458;
  wire n10460;
  wire n10461;
  wire [2:0] n10462;
  reg n10463;
  wire [31:0] n10464;
  wire n10466;
  wire [31:0] n10467;
  wire n10469;
  wire n10470;
  wire [30:0] n10471;
  wire [31:0] n10472;
  wire [31:0] n10473;
  wire n10474;
  wire [14:0] n10476;
  wire [14:0] n10477;
  wire [30:0] n10478;
  wire [63:0] n10479;
  wire n10480;
  wire [63:0] n10482;
  wire [63:0] n10484;
  wire [14:0] n10486;
  wire [63:0] n10487;
  wire n10489;
  wire [14:0] n10490;
  wire [63:0] n10491;
  wire n10492;
  wire n10493;
  wire [14:0] n10495;
  wire [63:0] n10497;
  wire n10499;
  wire n10500;
  wire [14:0] n10501;
  wire [63:0] n10502;
  wire n10503;
  wire n10505;
  wire n10506;
  wire n10507;
  wire n10508;
  wire n10509;
  wire n10511;
  wire n10513;
  wire n10515;
  wire n10516;
  wire n10517;
  wire n10518;
  wire [61:0] n10519;
  wire n10521;
  wire n10524;
  wire n10526;
  wire n10527;
  wire n10528;
  wire n10529;
  wire n10532;
  wire n10535;
  wire n10537;
  wire n10539;
  wire n10540;
  wire n10541;
  wire n10544;
  wire n10547;
  wire n10549;
  wire n10551;
  wire n10553;
  wire n10554;
  wire n10556;
  wire n10557;
  wire n10559;
  wire n10560;
  wire n10561;
  wire [61:0] n10562;
  wire n10564;
  wire n10567;
  wire n10571;
  wire n10573;
  wire n10575;
  wire n10577;
  wire n10579;
  wire n10580;
  wire n10583;
  wire n10586;
  wire n10589;
  wire [5:0] n10590;
  reg n10592;
  reg n10594;
  reg n10597;
  wire n10600;
  wire n10601;
  wire n10602;
  wire n10603;
  wire n10605;
  wire n10607;
  wire [14:0] n10609;
  wire [14:0] n10611;
  wire [63:0] n10614;
  wire n10616;
  wire [63:0] n10618;
  wire [14:0] n10619;
  wire [63:0] n10620;
  wire n10621;
  wire n10622;
  wire [63:0] n10623;
  wire n10624;
  wire n10626;
  wire n10628;
  wire n10629;
  wire n10630;
  wire n10631;
  wire n10632;
  wire n10634;
  wire n10636;
  wire [14:0] n10638;
  wire [14:0] n10640;
  wire [63:0] n10643;
  wire n10645;
  wire [63:0] n10647;
  wire [14:0] n10648;
  wire [63:0] n10649;
  wire n10650;
  wire n10651;
  wire [63:0] n10652;
  wire n10653;
  wire n10655;
  wire n10656;
  wire n10657;
  wire n10658;
  wire n10660;
  wire n10662;
  wire [14:0] n10664;
  wire [14:0] n10666;
  wire [63:0] n10669;
  wire n10671;
  wire [63:0] n10673;
  wire [14:0] n10674;
  wire [63:0] n10675;
  wire n10676;
  wire n10677;
  wire [63:0] n10678;
  wire n10679;
  wire n10681;
  wire [3:0] n10682;
  reg [14:0] n10683;
  reg [63:0] n10684;
  reg n10685;
  wire n10686;
  wire [14:0] n10688;
  wire [63:0] n10690;
  wire n10691;
  wire n10692;
  wire n10693;
  wire n10695;
  wire n10697;
  wire n10699;
  wire [14:0] n10701;
  wire [63:0] n10703;
  wire n10704;
  wire n10705;
  wire n10706;
  wire n10709;
  wire n10710;
  wire n10712;
  wire [14:0] n10714;
  wire [63:0] n10716;
  wire n10717;
  wire n10718;
  wire n10719;
  wire n10721;
  wire n10722;
  wire n10725;
  wire [15:0] n10726;
  wire [79:0] n10727;
  wire n10729;
  wire [5:0] n10730;
  reg [79:0] n10732;
  reg n10736;
  reg n10739;
  reg n10743;
  reg n10745;
  reg n10747;
  reg n10749;
  reg [14:0] n10751;
  reg [14:0] n10753;
  reg [14:0] n10755;
  reg [63:0] n10757;
  reg [63:0] n10759;
  reg [63:0] n10761;
  reg [2:0] n10767;
  reg [64:0] n10769;
  reg [64:0] n10775;
  reg [64:0] n10777;
  reg [14:0] n10779;
  reg n10783;
  reg n10785;
  reg n10787;
  reg [127:0] n10791;
  reg [7:0] n10793;
  reg n10796;
  reg n10799;
  reg n10802;
  reg n10805;
  reg n10808;
  wire n10943;
  wire n10944;
  wire n10945;
  reg n10946;
  wire n10947;
  wire n10948;
  wire n10949;
  reg n10950;
  wire n10951;
  wire n10952;
  wire n10953;
  reg n10954;
  wire n10955;
  wire n10956;
  wire [14:0] n10957;
  reg [14:0] n10958;
  wire n10959;
  wire n10960;
  wire [14:0] n10961;
  reg [14:0] n10962;
  wire n10963;
  wire n10964;
  wire [14:0] n10965;
  reg [14:0] n10966;
  wire n10967;
  wire n10968;
  wire [63:0] n10969;
  reg [63:0] n10970;
  wire n10971;
  wire n10972;
  wire [63:0] n10973;
  reg [63:0] n10974;
  wire n10975;
  wire n10976;
  wire [63:0] n10977;
  reg [63:0] n10978;
  wire [2:0] n10979;
  reg [2:0] n10980;
  wire n10982;
  wire n10983;
  wire [64:0] n10984;
  reg [64:0] n10985;
  wire n10995;
  wire n10996;
  wire [64:0] n10997;
  reg [64:0] n10998;
  wire n10999;
  wire n11000;
  wire [64:0] n11001;
  reg [64:0] n11002;
  wire n11003;
  wire n11004;
  wire [14:0] n11005;
  reg [14:0] n11006;
  wire n11011;
  wire n11012;
  wire n11013;
  reg n11014;
  wire n11015;
  wire n11016;
  wire n11017;
  reg n11018;
  wire n11019;
  wire n11020;
  wire n11021;
  reg n11022;
  wire n11029;
  wire n11030;
  wire [127:0] n11031;
  reg [127:0] n11032;
  wire n11039;
  wire n11040;
  wire [7:0] n11041;
  reg [7:0] n11042;
  wire n11043;
  reg n11044;
  wire n11045;
  reg n11046;
  wire n11047;
  reg n11048;
  wire n11049;
  reg n11050;
  wire n11051;
  reg n11052;
  wire [79:0] n11053;
  reg [79:0] n11054;
  wire n11055;
  reg n11056;
  wire n11057;
  reg n11058;
  wire n11059;
  reg n11060;
  assign result = n11054; //(module output)
  assign result_valid = n11056; //(module output)
  assign overflow = flags_overflow; //(module output)
  assign underflow = flags_underflow; //(module output)
  assign inexact = flags_inexact; //(module output)
  assign invalid = flags_invalid; //(module output)
  assign divide_by_zero = flags_div_by_zero; //(module output)
  assign quotient_byte = fmod_quotient; //(module output)
  assign operation_busy = n11058; //(module output)
  assign operation_done = n11060; //(module output)
  /* TG68K_FPU_ALU.vhd:1279:65  */
  assign sign_a = n10946; // (signal)
  /* TG68K_FPU_ALU.vhd:92:24  */
  assign sign_b = n10950; // (signal)
  /* TG68K_FPU_ALU.vhd:92:32  */
  assign sign_result = n10954; // (signal)
  /* TG68K_FPU_ALU.vhd:956:73  */
  assign exp_a = n10958; // (signal)
  /* TG68K_FPU_ALU.vhd:1105:81  */
  assign exp_b = n10962; // (signal)
  /* TG68K_FPU_ALU.vhd:93:30  */
  assign exp_result = n10966; // (signal)
  /* TG68K_FPU_ALU.vhd:94:16  */
  assign mant_a = n10970; // (signal)
  /* TG68K_FPU_ALU.vhd:94:24  */
  assign mant_b = n10974; // (signal)
  /* TG68K_FPU_ALU.vhd:94:32  */
  assign mant_result = n10978; // (signal)
  /* TG68K_FPU_ALU.vhd:105:16  */
  always @*
    alu_state = n10980; // (isignal)
  initial
    alu_state = 3'b000;
  /* TG68K_FPU_ALU.vhd:109:16  */
  assign mant_sum = n10985; // (signal)
  /* TG68K_FPU_ALU.vhd:115:16  */
  assign mant_a_aligned = n10998; // (signal)
  /* TG68K_FPU_ALU.vhd:115:32  */
  assign mant_b_aligned = n11002; // (signal)
  /* TG68K_FPU_ALU.vhd:116:16  */
  assign exp_larger = n11006; // (signal)
  /* TG68K_FPU_ALU.vhd:120:16  */
  assign guard_bit = n11014; // (signal)
  /* TG68K_FPU_ALU.vhd:120:27  */
  assign round_bit = n11018; // (signal)
  /* TG68K_FPU_ALU.vhd:120:38  */
  assign sticky_bit = n11022; // (signal)
  /* TG68K_FPU_ALU.vhd:127:16  */
  assign mult_result = n11032; // (signal)
  /* TG68K_FPU_ALU.vhd:138:16  */
  always @*
    fmod_quotient = n11042; // (isignal)
  initial
    fmod_quotient = 8'b00000000;
  /* TG68K_FPU_ALU.vhd:146:16  */
  assign is_zero_a = n7405; // (signal)
  /* TG68K_FPU_ALU.vhd:146:27  */
  assign is_zero_b = n7465; // (signal)
  /* TG68K_FPU_ALU.vhd:147:16  */
  assign is_inf_a = n7407; // (signal)
  /* TG68K_FPU_ALU.vhd:147:26  */
  assign is_inf_b = n7467; // (signal)
  /* TG68K_FPU_ALU.vhd:148:16  */
  assign is_nan_a = n7409; // (signal)
  /* TG68K_FPU_ALU.vhd:148:26  */
  assign is_nan_b = n7469; // (signal)
  /* TG68K_FPU_ALU.vhd:149:16  */
  assign is_denorm_a = n7411; // (signal)
  /* TG68K_FPU_ALU.vhd:149:29  */
  assign is_denorm_b = n7471; // (signal)
  /* TG68K_FPU_ALU.vhd:150:16  */
  assign is_snan_a = n7413; // (signal)
  /* TG68K_FPU_ALU.vhd:150:27  */
  assign is_snan_b = n7473; // (signal)
  /* TG68K_FPU_ALU.vhd:159:16  */
  assign flags_overflow = n11044; // (signal)
  /* TG68K_FPU_ALU.vhd:160:16  */
  assign flags_underflow = n11046; // (signal)
  /* TG68K_FPU_ALU.vhd:161:16  */
  assign flags_inexact = n11048; // (signal)
  /* TG68K_FPU_ALU.vhd:162:16  */
  assign flags_invalid = n11050; // (signal)
  /* TG68K_FPU_ALU.vhd:163:16  */
  assign flags_div_by_zero = n11052; // (signal)
  /* TG68K_FPU_ALU.vhd:171:29  */
  assign n7356 = operand_a[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:171:44  */
  assign n7358 = n7356 == 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:172:37  */
  assign n7359 = operand_a[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:172:51  */
  assign n7361 = n7359 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:172:25  */
  assign n7364 = n7361 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:172:25  */
  assign n7367 = n7361 ? 1'b0 : 1'b1;
  /* TG68K_FPU_ALU.vhd:183:32  */
  assign n7368 = operand_a[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:183:47  */
  assign n7370 = n7368 == 15'b111111111111111;
  /* TG68K_FPU_ALU.vhd:186:37  */
  assign n7371 = operand_a[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:186:51  */
  assign n7373 = n7371 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:197:45  */
  assign n7374 = operand_a[62]; // extract
  /* TG68K_FPU_ALU.vhd:197:50  */
  assign n7375 = ~n7374;
  /* TG68K_FPU_ALU.vhd:197:69  */
  assign n7376 = operand_a[61:0]; // extract
  /* TG68K_FPU_ALU.vhd:197:83  */
  assign n7378 = n7376 != 62'b00000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:197:56  */
  assign n7379 = n7378 & n7375;
  /* TG68K_FPU_ALU.vhd:197:33  */
  assign n7382 = n7379 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:186:25  */
  assign n7388 = n7373 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:186:25  */
  assign n7391 = n7373 ? 1'b0 : 1'b1;
  /* TG68K_FPU_ALU.vhd:186:25  */
  assign n7393 = n7373 ? 1'b0 : n7382;
  /* TG68K_FPU_ALU.vhd:183:17  */
  assign n7397 = n7370 ? n7388 : 1'b0;
  /* TG68K_FPU_ALU.vhd:183:17  */
  assign n7399 = n7370 ? n7391 : 1'b0;
  /* TG68K_FPU_ALU.vhd:183:17  */
  assign n7401 = n7370 ? n7393 : 1'b0;
  /* TG68K_FPU_ALU.vhd:171:17  */
  assign n7405 = n7358 ? n7364 : 1'b0;
  /* TG68K_FPU_ALU.vhd:171:17  */
  assign n7407 = n7358 ? 1'b0 : n7397;
  /* TG68K_FPU_ALU.vhd:171:17  */
  assign n7409 = n7358 ? 1'b0 : n7399;
  /* TG68K_FPU_ALU.vhd:171:17  */
  assign n7411 = n7358 ? n7367 : 1'b0;
  /* TG68K_FPU_ALU.vhd:171:17  */
  assign n7413 = n7358 ? 1'b0 : n7401;
  /* TG68K_FPU_ALU.vhd:215:29  */
  assign n7416 = operand_b[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:215:44  */
  assign n7418 = n7416 == 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:216:37  */
  assign n7419 = operand_b[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:216:51  */
  assign n7421 = n7419 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:216:25  */
  assign n7424 = n7421 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:216:25  */
  assign n7427 = n7421 ? 1'b0 : 1'b1;
  /* TG68K_FPU_ALU.vhd:227:32  */
  assign n7428 = operand_b[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:227:47  */
  assign n7430 = n7428 == 15'b111111111111111;
  /* TG68K_FPU_ALU.vhd:230:37  */
  assign n7431 = operand_b[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:230:51  */
  assign n7433 = n7431 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:241:45  */
  assign n7434 = operand_b[62]; // extract
  /* TG68K_FPU_ALU.vhd:241:50  */
  assign n7435 = ~n7434;
  /* TG68K_FPU_ALU.vhd:241:69  */
  assign n7436 = operand_b[61:0]; // extract
  /* TG68K_FPU_ALU.vhd:241:83  */
  assign n7438 = n7436 != 62'b00000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:241:56  */
  assign n7439 = n7438 & n7435;
  /* TG68K_FPU_ALU.vhd:241:33  */
  assign n7442 = n7439 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:230:25  */
  assign n7448 = n7433 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:230:25  */
  assign n7451 = n7433 ? 1'b0 : 1'b1;
  /* TG68K_FPU_ALU.vhd:230:25  */
  assign n7453 = n7433 ? 1'b0 : n7442;
  /* TG68K_FPU_ALU.vhd:227:17  */
  assign n7457 = n7430 ? n7448 : 1'b0;
  /* TG68K_FPU_ALU.vhd:227:17  */
  assign n7459 = n7430 ? n7451 : 1'b0;
  /* TG68K_FPU_ALU.vhd:227:17  */
  assign n7461 = n7430 ? n7453 : 1'b0;
  /* TG68K_FPU_ALU.vhd:215:17  */
  assign n7465 = n7418 ? n7424 : 1'b0;
  /* TG68K_FPU_ALU.vhd:215:17  */
  assign n7467 = n7418 ? 1'b0 : n7457;
  /* TG68K_FPU_ALU.vhd:215:17  */
  assign n7469 = n7418 ? 1'b0 : n7459;
  /* TG68K_FPU_ALU.vhd:215:17  */
  assign n7471 = n7418 ? n7427 : 1'b0;
  /* TG68K_FPU_ALU.vhd:215:17  */
  assign n7473 = n7418 ? 1'b0 : n7461;
  /* TG68K_FPU_ALU.vhd:267:27  */
  assign n7481 = ~nreset;
  /* TG68K_FPU_ALU.vhd:289:49  */
  assign n7485 = start_operation ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:289:49  */
  assign n7488 = start_operation ? 3'b001 : alu_state;
  /* TG68K_FPU_ALU.vhd:284:41  */
  assign n7490 = alu_state == 3'b000;
  /* TG68K_FPU_ALU.vhd:294:41  */
  assign n7492 = alu_state == 3'b001;
  /* TG68K_FPU_ALU.vhd:307:68  */
  assign n7493 = operand_a[79]; // extract
  /* TG68K_FPU_ALU.vhd:308:67  */
  assign n7494 = operand_a[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:309:68  */
  assign n7495 = operand_a[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:311:68  */
  assign n7496 = operand_b[79]; // extract
  /* TG68K_FPU_ALU.vhd:312:67  */
  assign n7497 = operand_b[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:313:68  */
  assign n7498 = operand_b[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:316:67  */
  assign n7500 = operation_code == 7'b0000000;
  /* TG68K_FPU_ALU.vhd:318:81  */
  assign n7501 = operand_a[79]; // extract
  /* TG68K_FPU_ALU.vhd:319:80  */
  assign n7502 = operand_a[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:320:81  */
  assign n7503 = operand_a[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:322:70  */
  assign n7505 = operation_code == 7'b0100010;
  /* TG68K_FPU_ALU.vhd:322:80  */
  assign n7506 = is_zero_b & n7505;
  /* TG68K_FPU_ALU.vhd:322:116  */
  assign n7507 = ~is_denorm_a;
  /* TG68K_FPU_ALU.vhd:322:100  */
  assign n7508 = n7507 & n7506;
  /* TG68K_FPU_ALU.vhd:324:81  */
  assign n7509 = operand_a[79]; // extract
  /* TG68K_FPU_ALU.vhd:325:80  */
  assign n7510 = operand_a[78:64]; // extract
  /* TG68K_FPU_ALU.vhd:326:81  */
  assign n7511 = operand_a[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:328:70  */
  assign n7513 = operation_code == 7'b0100011;
  /* TG68K_FPU_ALU.vhd:328:101  */
  assign n7514 = is_zero_a | is_zero_b;
  /* TG68K_FPU_ALU.vhd:328:80  */
  assign n7515 = n7514 & n7513;
  /* TG68K_FPU_ALU.vhd:330:81  */
  assign n7516 = operand_a[79]; // extract
  /* TG68K_FPU_ALU.vhd:330:99  */
  assign n7517 = operand_b[79]; // extract
  /* TG68K_FPU_ALU.vhd:330:86  */
  assign n7518 = n7516 ^ n7517;
  /* TG68K_FPU_ALU.vhd:328:49  */
  assign n7519 = n7515 ? n7518 : sign_result;
  /* TG68K_FPU_ALU.vhd:328:49  */
  assign n7521 = n7515 ? 15'b000000000000000 : exp_result;
  /* TG68K_FPU_ALU.vhd:328:49  */
  assign n7523 = n7515 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : mant_result;
  /* TG68K_FPU_ALU.vhd:328:49  */
  assign n7526 = n7515 ? 3'b100 : 3'b011;
  /* TG68K_FPU_ALU.vhd:322:49  */
  assign n7527 = n7508 ? n7509 : n7519;
  /* TG68K_FPU_ALU.vhd:322:49  */
  assign n7528 = n7508 ? n7510 : n7521;
  /* TG68K_FPU_ALU.vhd:322:49  */
  assign n7529 = n7508 ? n7511 : n7523;
  /* TG68K_FPU_ALU.vhd:322:49  */
  assign n7531 = n7508 ? 3'b100 : n7526;
  /* TG68K_FPU_ALU.vhd:316:49  */
  assign n7532 = n7500 ? n7501 : n7527;
  /* TG68K_FPU_ALU.vhd:316:49  */
  assign n7533 = n7500 ? n7502 : n7528;
  /* TG68K_FPU_ALU.vhd:316:49  */
  assign n7534 = n7500 ? n7503 : n7529;
  /* TG68K_FPU_ALU.vhd:316:49  */
  assign n7536 = n7500 ? 3'b100 : n7531;
  /* TG68K_FPU_ALU.vhd:304:41  */
  assign n7538 = alu_state == 3'b010;
  /* TG68K_FPU_ALU.vhd:340:57  */
  assign n7540 = operation_code == 7'b0000000;
  /* TG68K_FPU_ALU.vhd:347:57  */
  assign n7542 = operation_code == 7'b0011000;
  /* TG68K_FPU_ALU.vhd:356:80  */
  assign n7543 = ~sign_a;
  /* TG68K_FPU_ALU.vhd:354:57  */
  assign n7545 = operation_code == 7'b0011010;
  /* TG68K_FPU_ALU.vhd:363:85  */
  assign n7546 = ~is_zero_a;
  /* TG68K_FPU_ALU.vhd:363:81  */
  assign n7547 = n7546 & sign_a;
  /* TG68K_FPU_ALU.vhd:385:85  */
  assign n7548 = {16'b0, exp_a};  //  uext
  /* TG68K_FPU_ALU.vhd:385:113  */
  assign n7549 = {1'b0, n7548};  //  uext
  /* TG68K_FPU_ALU.vhd:385:113  */
  assign n7551 = n7549 - 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:386:125  */
  assign n7553 = $signed(n7551) / $signed(32'b00000000000000000000000000000010); // sdiv
  /* TG68K_FPU_ALU.vhd:386:129  */
  assign n7555 = n7553 + 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:386:116  */
  assign n7556 = n7555[30:0];  // trunc
  /* TG68K_FPU_ALU.vhd:386:104  */
  assign n7557 = n7556[14:0];  // trunc
  /* TG68K_FPU_ALU.vhd:390:82  */
  assign n7558 = mant_a[63:62]; // extract
  /* TG68K_FPU_ALU.vhd:390:97  */
  assign n7560 = n7558 == 2'b11;
  /* TG68K_FPU_ALU.vhd:393:85  */
  assign n7561 = mant_a[63:62]; // extract
  /* TG68K_FPU_ALU.vhd:393:100  */
  assign n7563 = n7561 == 2'b10;
  /* TG68K_FPU_ALU.vhd:396:85  */
  assign n7564 = mant_a[63:62]; // extract
  /* TG68K_FPU_ALU.vhd:396:100  */
  assign n7566 = n7564 == 2'b01;
  /* TG68K_FPU_ALU.vhd:396:73  */
  assign n7569 = n7566 ? 64'b1000111101011100001010001111010111000010100011110101110000101001 : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:393:73  */
  assign n7571 = n7563 ? 64'b1001110110001001110110001001110110001001110110001001110110001010 : n7569;
  /* TG68K_FPU_ALU.vhd:390:73  */
  assign n7573 = n7560 ? 64'b1010100011110101110000101000111101011100001010001111010111000011 : n7571;
  /* TG68K_FPU_ALU.vhd:405:81  */
  assign n7574 = exp_a[0]; // extract
  /* TG68K_FPU_ALU.vhd:408:157  */
  assign n7575 = mant_result[63:1]; // extract
  /* TG68K_FPU_ALU.vhd:408:135  */
  assign n7576 = {1'b0, n7575};  //  uext
  /* TG68K_FPU_ALU.vhd:408:135  */
  assign n7577 = mant_result + n7576;
  /* TG68K_FPU_ALU.vhd:405:73  */
  assign n7578 = n7574 ? n7577 : n7573;
  /* TG68K_FPU_ALU.vhd:374:65  */
  assign n7580 = is_inf_a ? 15'b111111111111111 : n7557;
  /* TG68K_FPU_ALU.vhd:374:65  */
  assign n7582 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7578;
  /* TG68K_FPU_ALU.vhd:374:65  */
  assign n7584 = is_inf_a ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:369:65  */
  assign n7587 = is_zero_a ? 15'b000000000000000 : n7580;
  /* TG68K_FPU_ALU.vhd:369:65  */
  assign n7589 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7582;
  /* TG68K_FPU_ALU.vhd:369:65  */
  assign n7590 = is_zero_a ? flags_inexact : n7584;
  /* TG68K_FPU_ALU.vhd:363:65  */
  assign n7593 = n7547 ? 15'b111111111111111 : n7587;
  /* TG68K_FPU_ALU.vhd:363:65  */
  assign n7595 = n7547 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n7589;
  /* TG68K_FPU_ALU.vhd:363:65  */
  assign n7596 = n7547 ? flags_inexact : n7590;
  /* TG68K_FPU_ALU.vhd:363:65  */
  assign n7598 = n7547 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:361:57  */
  assign n7601 = operation_code == 7'b0000100;
  /* TG68K_FPU_ALU.vhd:417:83  */
  assign n7602 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:420:92  */
  assign n7603 = is_snan_a | is_snan_b;
  /* TG68K_FPU_ALU.vhd:420:73  */
  assign n7605 = n7603 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:427:86  */
  assign n7606 = is_inf_b & is_inf_a;
  /* TG68K_FPU_ALU.vhd:429:83  */
  assign n7607 = sign_a == sign_b;
  /* TG68K_FPU_ALU.vhd:429:73  */
  assign n7609 = n7607 ? sign_a : 1'b0;
  /* TG68K_FPU_ALU.vhd:429:73  */
  assign n7612 = n7607 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:429:73  */
  assign n7614 = n7607 ? flags_invalid : 1'b1;
  /* TG68K_FPU_ALU.vhd:451:103  */
  assign n7615 = ~is_denorm_b;
  /* TG68K_FPU_ALU.vhd:451:87  */
  assign n7616 = n7615 & is_zero_a;
  /* TG68K_FPU_ALU.vhd:456:103  */
  assign n7617 = ~is_denorm_a;
  /* TG68K_FPU_ALU.vhd:456:87  */
  assign n7618 = n7617 & is_zero_b;
  /* TG68K_FPU_ALU.vhd:461:89  */
  assign n7619 = is_denorm_a | is_denorm_b;
  /* TG68K_FPU_ALU.vhd:465:82  */
  assign n7621 = exp_a == 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:467:103  */
  assign n7623 = {1'b0, mant_a};
  /* TG68K_FPU_ALU.vhd:469:103  */
  assign n7625 = {1'b1, mant_a};
  /* TG68K_FPU_ALU.vhd:465:73  */
  assign n7626 = n7621 ? n7623 : n7625;
  /* TG68K_FPU_ALU.vhd:471:82  */
  assign n7628 = exp_b == 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:473:103  */
  assign n7630 = {1'b0, mant_b};
  /* TG68K_FPU_ALU.vhd:475:103  */
  assign n7632 = {1'b1, mant_b};
  /* TG68K_FPU_ALU.vhd:471:73  */
  assign n7633 = n7628 ? n7630 : n7632;
  /* TG68K_FPU_ALU.vhd:480:83  */
  assign n7634 = sign_a == sign_b;
  /* TG68K_FPU_ALU.vhd:482:108  */
  assign n7635 = mant_a_aligned + mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:486:99  */
  assign n7636 = $unsigned(mant_a_aligned) >= $unsigned(mant_b_aligned);
  /* TG68K_FPU_ALU.vhd:487:116  */
  assign n7637 = mant_a_aligned - mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:490:116  */
  assign n7638 = mant_b_aligned - mant_a_aligned;
  /* TG68K_FPU_ALU.vhd:486:81  */
  assign n7639 = n7636 ? sign_a : sign_b;
  /* TG68K_FPU_ALU.vhd:486:81  */
  assign n7640 = n7636 ? n7637 : n7638;
  /* TG68K_FPU_ALU.vhd:480:73  */
  assign n7641 = n7634 ? sign_a : n7639;
  /* TG68K_FPU_ALU.vhd:480:73  */
  assign n7642 = n7634 ? n7635 : n7640;
  /* TG68K_FPU_ALU.vhd:498:82  */
  assign n7643 = $unsigned(exp_a) >= $unsigned(exp_b);
  /* TG68K_FPU_ALU.vhd:503:103  */
  assign n7646 = {1'b1, mant_a};
  /* TG68K_FPU_ALU.vhd:505:90  */
  assign n7647 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:505:98  */
  assign n7649 = $unsigned(n7647) > $unsigned(15'b000000000111111);
  /* TG68K_FPU_ALU.vhd:510:149  */
  assign n7654 = {1'b1, mant_b};
  /* TG68K_FPU_ALU.vhd:510:186  */
  assign n7655 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:510:160  */
  assign n7656 = {16'b0, n7655};  //  uext
  /* TG68K_FPU_ALU.vhd:510:124  */
  assign n7657 = n7654 >> n7656;
  /* TG68K_FPU_ALU.vhd:505:81  */
  assign n7660 = n7649 ? 65'b00000000000000000000000000000000000000000000000000000000000000000 : n7657;
  /* TG68K_FPU_ALU.vhd:517:103  */
  assign n7663 = {1'b1, mant_b};
  /* TG68K_FPU_ALU.vhd:519:90  */
  assign n7664 = exp_b - exp_a;
  /* TG68K_FPU_ALU.vhd:519:98  */
  assign n7666 = $unsigned(n7664) > $unsigned(15'b000000000111111);
  /* TG68K_FPU_ALU.vhd:524:149  */
  assign n7671 = {1'b1, mant_a};
  /* TG68K_FPU_ALU.vhd:524:186  */
  assign n7672 = exp_b - exp_a;
  /* TG68K_FPU_ALU.vhd:524:160  */
  assign n7673 = {16'b0, n7672};  //  uext
  /* TG68K_FPU_ALU.vhd:524:124  */
  assign n7674 = n7671 >> n7673;
  /* TG68K_FPU_ALU.vhd:519:81  */
  assign n7677 = n7666 ? 65'b00000000000000000000000000000000000000000000000000000000000000000 : n7674;
  /* TG68K_FPU_ALU.vhd:498:73  */
  assign n7680 = n7643 ? n7646 : n7677;
  /* TG68K_FPU_ALU.vhd:498:73  */
  assign n7681 = n7643 ? n7660 : n7663;
  /* TG68K_FPU_ALU.vhd:498:73  */
  assign n7682 = n7643 ? exp_a : exp_b;
  /* TG68K_FPU_ALU.vhd:529:84  */
  assign n7684 = sign_a == sign_b;
  /* TG68K_FPU_ALU.vhd:531:108  */
  assign n7685 = mant_a_aligned + mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:535:99  */
  assign n7686 = $unsigned(mant_a_aligned) >= $unsigned(mant_b_aligned);
  /* TG68K_FPU_ALU.vhd:536:116  */
  assign n7687 = mant_a_aligned - mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:539:116  */
  assign n7688 = mant_b_aligned - mant_a_aligned;
  /* TG68K_FPU_ALU.vhd:535:81  */
  assign n7689 = n7686 ? sign_a : sign_b;
  /* TG68K_FPU_ALU.vhd:535:81  */
  assign n7690 = n7686 ? n7687 : n7688;
  /* TG68K_FPU_ALU.vhd:529:73  */
  assign n7691 = n7684 ? sign_a : n7689;
  /* TG68K_FPU_ALU.vhd:529:73  */
  assign n7692 = n7684 ? n7685 : n7690;
  /* TG68K_FPU_ALU.vhd:545:84  */
  assign n7693 = mant_sum[64]; // extract
  /* TG68K_FPU_ALU.vhd:547:133  */
  assign n7695 = exp_larger + 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:548:104  */
  assign n7696 = mant_sum[64:1]; // extract
  /* TG68K_FPU_ALU.vhd:549:87  */
  assign n7697 = mant_sum[63]; // extract
  /* TG68K_FPU_ALU.vhd:549:92  */
  assign n7698 = ~n7697;
  /* TG68K_FPU_ALU.vhd:551:133  */
  assign n7700 = exp_larger - 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:552:104  */
  assign n7701 = mant_sum[62:0]; // extract
  /* TG68K_FPU_ALU.vhd:552:118  */
  assign n7703 = {n7701, 1'b0};
  /* TG68K_FPU_ALU.vhd:556:104  */
  assign n7704 = mant_sum[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:549:73  */
  assign n7705 = n7698 ? n7700 : exp_larger;
  /* TG68K_FPU_ALU.vhd:549:73  */
  assign n7706 = n7698 ? n7703 : n7704;
  /* TG68K_FPU_ALU.vhd:545:73  */
  assign n7707 = n7693 ? n7695 : n7705;
  /* TG68K_FPU_ALU.vhd:545:73  */
  assign n7708 = n7693 ? n7696 : n7706;
  /* TG68K_FPU_ALU.vhd:461:65  */
  assign n7709 = n7619 ? n7641 : n7691;
  /* TG68K_FPU_ALU.vhd:461:65  */
  assign n7710 = n7619 ? exp_larger : n7707;
  /* TG68K_FPU_ALU.vhd:461:65  */
  assign n7711 = n7619 ? mant_result : n7708;
  /* TG68K_FPU_ALU.vhd:461:65  */
  assign n7712 = n7619 ? n7642 : n7692;
  /* TG68K_FPU_ALU.vhd:461:65  */
  assign n7715 = n7619 ? n7626 : n7680;
  /* TG68K_FPU_ALU.vhd:461:65  */
  assign n7716 = n7619 ? n7633 : n7681;
  /* TG68K_FPU_ALU.vhd:461:65  */
  assign n7718 = n7619 ? 15'b000000000000001 : n7682;
  /* TG68K_FPU_ALU.vhd:456:65  */
  assign n7720 = n7618 ? sign_a : n7709;
  /* TG68K_FPU_ALU.vhd:456:65  */
  assign n7721 = n7618 ? exp_a : n7710;
  /* TG68K_FPU_ALU.vhd:456:65  */
  assign n7722 = n7618 ? mant_a : n7711;
  /* TG68K_FPU_ALU.vhd:456:65  */
  assign n7723 = n7618 ? mant_sum : n7712;
  /* TG68K_FPU_ALU.vhd:456:65  */
  assign n7726 = n7618 ? mant_a_aligned : n7715;
  /* TG68K_FPU_ALU.vhd:456:65  */
  assign n7727 = n7618 ? mant_b_aligned : n7716;
  /* TG68K_FPU_ALU.vhd:456:65  */
  assign n7728 = n7618 ? exp_larger : n7718;
  /* TG68K_FPU_ALU.vhd:451:65  */
  assign n7730 = n7616 ? sign_b : n7720;
  /* TG68K_FPU_ALU.vhd:451:65  */
  assign n7731 = n7616 ? exp_b : n7721;
  /* TG68K_FPU_ALU.vhd:451:65  */
  assign n7732 = n7616 ? mant_b : n7722;
  /* TG68K_FPU_ALU.vhd:451:65  */
  assign n7733 = n7616 ? mant_sum : n7723;
  /* TG68K_FPU_ALU.vhd:451:65  */
  assign n7736 = n7616 ? mant_a_aligned : n7726;
  /* TG68K_FPU_ALU.vhd:451:65  */
  assign n7737 = n7616 ? mant_b_aligned : n7727;
  /* TG68K_FPU_ALU.vhd:451:65  */
  assign n7738 = n7616 ? exp_larger : n7728;
  /* TG68K_FPU_ALU.vhd:446:65  */
  assign n7740 = is_inf_b ? sign_b : n7730;
  /* TG68K_FPU_ALU.vhd:446:65  */
  assign n7742 = is_inf_b ? 15'b111111111111111 : n7731;
  /* TG68K_FPU_ALU.vhd:446:65  */
  assign n7744 = is_inf_b ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7732;
  /* TG68K_FPU_ALU.vhd:446:65  */
  assign n7745 = is_inf_b ? mant_sum : n7733;
  /* TG68K_FPU_ALU.vhd:446:65  */
  assign n7748 = is_inf_b ? mant_a_aligned : n7736;
  /* TG68K_FPU_ALU.vhd:446:65  */
  assign n7749 = is_inf_b ? mant_b_aligned : n7737;
  /* TG68K_FPU_ALU.vhd:446:65  */
  assign n7750 = is_inf_b ? exp_larger : n7738;
  /* TG68K_FPU_ALU.vhd:441:65  */
  assign n7752 = is_inf_a ? sign_a : n7740;
  /* TG68K_FPU_ALU.vhd:441:65  */
  assign n7754 = is_inf_a ? 15'b111111111111111 : n7742;
  /* TG68K_FPU_ALU.vhd:441:65  */
  assign n7756 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7744;
  /* TG68K_FPU_ALU.vhd:441:65  */
  assign n7757 = is_inf_a ? mant_sum : n7745;
  /* TG68K_FPU_ALU.vhd:441:65  */
  assign n7760 = is_inf_a ? mant_a_aligned : n7748;
  /* TG68K_FPU_ALU.vhd:441:65  */
  assign n7761 = is_inf_a ? mant_b_aligned : n7749;
  /* TG68K_FPU_ALU.vhd:441:65  */
  assign n7762 = is_inf_a ? exp_larger : n7750;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7764 = n7606 ? n7609 : n7752;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7766 = n7606 ? 15'b111111111111111 : n7754;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7767 = n7606 ? n7612 : n7756;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7768 = n7606 ? mant_sum : n7757;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7771 = n7606 ? mant_a_aligned : n7760;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7772 = n7606 ? mant_b_aligned : n7761;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7773 = n7606 ? exp_larger : n7762;
  /* TG68K_FPU_ALU.vhd:427:65  */
  assign n7775 = n7606 ? n7614 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7777 = n7602 ? 1'b0 : n7764;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7779 = n7602 ? 15'b111111111111111 : n7766;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7781 = n7602 ? 64'b1100000000000000000000000000000000000000000000000000000000000000 : n7767;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7782 = n7602 ? mant_sum : n7768;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7785 = n7602 ? mant_a_aligned : n7771;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7786 = n7602 ? mant_b_aligned : n7772;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7787 = n7602 ? exp_larger : n7773;
  /* TG68K_FPU_ALU.vhd:417:65  */
  assign n7789 = n7602 ? n7605 : n7775;
  /* TG68K_FPU_ALU.vhd:415:57  */
  assign n7791 = operation_code == 7'b0100010;
  /* TG68K_FPU_ALU.vhd:563:83  */
  assign n7792 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:569:86  */
  assign n7793 = is_inf_b & is_inf_a;
  /* TG68K_FPU_ALU.vhd:571:83  */
  assign n7794 = sign_a == sign_b;
  /* TG68K_FPU_ALU.vhd:571:73  */
  assign n7796 = n7794 ? 1'b0 : sign_a;
  /* TG68K_FPU_ALU.vhd:571:73  */
  assign n7799 = n7794 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7801 = n7944 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:590:88  */
  assign n7802 = ~sign_b;
  /* TG68K_FPU_ALU.vhd:593:103  */
  assign n7803 = ~is_denorm_b;
  /* TG68K_FPU_ALU.vhd:593:87  */
  assign n7804 = n7803 & is_zero_a;
  /* TG68K_FPU_ALU.vhd:595:88  */
  assign n7805 = ~sign_b;
  /* TG68K_FPU_ALU.vhd:598:103  */
  assign n7806 = ~is_denorm_a;
  /* TG68K_FPU_ALU.vhd:598:87  */
  assign n7807 = n7806 & is_zero_b;
  /* TG68K_FPU_ALU.vhd:603:89  */
  assign n7808 = is_denorm_a | is_denorm_b;
  /* TG68K_FPU_ALU.vhd:607:82  */
  assign n7810 = exp_a == 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:609:103  */
  assign n7812 = {1'b0, mant_a};
  /* TG68K_FPU_ALU.vhd:611:103  */
  assign n7814 = {1'b1, mant_a};
  /* TG68K_FPU_ALU.vhd:607:73  */
  assign n7815 = n7810 ? n7812 : n7814;
  /* TG68K_FPU_ALU.vhd:613:82  */
  assign n7817 = exp_b == 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:615:103  */
  assign n7819 = {1'b0, mant_b};
  /* TG68K_FPU_ALU.vhd:617:103  */
  assign n7821 = {1'b1, mant_b};
  /* TG68K_FPU_ALU.vhd:613:73  */
  assign n7822 = n7817 ? n7819 : n7821;
  /* TG68K_FPU_ALU.vhd:622:83  */
  assign n7823 = sign_a == sign_b;
  /* TG68K_FPU_ALU.vhd:624:99  */
  assign n7824 = $unsigned(mant_a_aligned) >= $unsigned(mant_b_aligned);
  /* TG68K_FPU_ALU.vhd:625:116  */
  assign n7825 = mant_a_aligned - mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:628:116  */
  assign n7826 = mant_b_aligned - mant_a_aligned;
  /* TG68K_FPU_ALU.vhd:629:104  */
  assign n7827 = ~sign_a;
  /* TG68K_FPU_ALU.vhd:624:81  */
  assign n7828 = n7824 ? sign_a : n7827;
  /* TG68K_FPU_ALU.vhd:624:81  */
  assign n7829 = n7824 ? n7825 : n7826;
  /* TG68K_FPU_ALU.vhd:633:108  */
  assign n7830 = mant_a_aligned + mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:622:73  */
  assign n7831 = n7823 ? n7828 : sign_a;
  /* TG68K_FPU_ALU.vhd:622:73  */
  assign n7832 = n7823 ? n7829 : n7830;
  /* TG68K_FPU_ALU.vhd:640:82  */
  assign n7833 = $unsigned(exp_a) >= $unsigned(exp_b);
  /* TG68K_FPU_ALU.vhd:644:103  */
  assign n7836 = {1'b1, mant_a};
  /* TG68K_FPU_ALU.vhd:646:90  */
  assign n7837 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:646:98  */
  assign n7839 = $unsigned(n7837) > $unsigned(15'b000000000111111);
  /* TG68K_FPU_ALU.vhd:649:149  */
  assign n7841 = {1'b1, mant_b};
  /* TG68K_FPU_ALU.vhd:649:186  */
  assign n7842 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:649:160  */
  assign n7843 = {16'b0, n7842};  //  uext
  /* TG68K_FPU_ALU.vhd:649:124  */
  assign n7844 = n7841 >> n7843;
  /* TG68K_FPU_ALU.vhd:646:81  */
  assign n7846 = n7839 ? 65'b00000000000000000000000000000000000000000000000000000000000000000 : n7844;
  /* TG68K_FPU_ALU.vhd:655:103  */
  assign n7849 = {1'b1, mant_b};
  /* TG68K_FPU_ALU.vhd:657:90  */
  assign n7850 = exp_b - exp_a;
  /* TG68K_FPU_ALU.vhd:657:98  */
  assign n7852 = $unsigned(n7850) > $unsigned(15'b000000000111111);
  /* TG68K_FPU_ALU.vhd:660:149  */
  assign n7854 = {1'b1, mant_a};
  /* TG68K_FPU_ALU.vhd:660:186  */
  assign n7855 = exp_b - exp_a;
  /* TG68K_FPU_ALU.vhd:660:160  */
  assign n7856 = {16'b0, n7855};  //  uext
  /* TG68K_FPU_ALU.vhd:660:124  */
  assign n7857 = n7854 >> n7856;
  /* TG68K_FPU_ALU.vhd:657:81  */
  assign n7859 = n7852 ? 65'b00000000000000000000000000000000000000000000000000000000000000000 : n7857;
  /* TG68K_FPU_ALU.vhd:640:73  */
  assign n7861 = n7833 ? n7836 : n7859;
  /* TG68K_FPU_ALU.vhd:640:73  */
  assign n7862 = n7833 ? n7846 : n7849;
  /* TG68K_FPU_ALU.vhd:640:73  */
  assign n7863 = n7833 ? exp_a : exp_b;
  /* TG68K_FPU_ALU.vhd:665:84  */
  assign n7864 = sign_a != sign_b;
  /* TG68K_FPU_ALU.vhd:667:108  */
  assign n7865 = mant_a_aligned + mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:671:99  */
  assign n7866 = $unsigned(mant_a_aligned) >= $unsigned(mant_b_aligned);
  /* TG68K_FPU_ALU.vhd:672:116  */
  assign n7867 = mant_a_aligned - mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:675:116  */
  assign n7868 = mant_b_aligned - mant_a_aligned;
  /* TG68K_FPU_ALU.vhd:676:104  */
  assign n7869 = ~sign_a;
  /* TG68K_FPU_ALU.vhd:671:81  */
  assign n7870 = n7866 ? sign_a : n7869;
  /* TG68K_FPU_ALU.vhd:671:81  */
  assign n7871 = n7866 ? n7867 : n7868;
  /* TG68K_FPU_ALU.vhd:665:73  */
  assign n7872 = n7864 ? sign_a : n7870;
  /* TG68K_FPU_ALU.vhd:665:73  */
  assign n7873 = n7864 ? n7865 : n7871;
  /* TG68K_FPU_ALU.vhd:681:84  */
  assign n7874 = mant_sum[64]; // extract
  /* TG68K_FPU_ALU.vhd:683:133  */
  assign n7876 = exp_larger + 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:684:104  */
  assign n7877 = mant_sum[64:1]; // extract
  /* TG68K_FPU_ALU.vhd:685:87  */
  assign n7878 = mant_sum[63]; // extract
  /* TG68K_FPU_ALU.vhd:685:92  */
  assign n7879 = ~n7878;
  /* TG68K_FPU_ALU.vhd:687:133  */
  assign n7881 = exp_larger - 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:688:104  */
  assign n7882 = mant_sum[62:0]; // extract
  /* TG68K_FPU_ALU.vhd:688:118  */
  assign n7884 = {n7882, 1'b0};
  /* TG68K_FPU_ALU.vhd:692:104  */
  assign n7885 = mant_sum[63:0]; // extract
  /* TG68K_FPU_ALU.vhd:685:73  */
  assign n7886 = n7879 ? n7881 : exp_larger;
  /* TG68K_FPU_ALU.vhd:685:73  */
  assign n7887 = n7879 ? n7884 : n7885;
  /* TG68K_FPU_ALU.vhd:681:73  */
  assign n7888 = n7874 ? n7876 : n7886;
  /* TG68K_FPU_ALU.vhd:681:73  */
  assign n7889 = n7874 ? n7877 : n7887;
  /* TG68K_FPU_ALU.vhd:603:65  */
  assign n7890 = n7808 ? n7831 : n7872;
  /* TG68K_FPU_ALU.vhd:603:65  */
  assign n7891 = n7808 ? exp_larger : n7888;
  /* TG68K_FPU_ALU.vhd:603:65  */
  assign n7892 = n7808 ? mant_result : n7889;
  /* TG68K_FPU_ALU.vhd:603:65  */
  assign n7893 = n7808 ? n7832 : n7873;
  /* TG68K_FPU_ALU.vhd:603:65  */
  assign n7895 = n7808 ? n7815 : n7861;
  /* TG68K_FPU_ALU.vhd:603:65  */
  assign n7896 = n7808 ? n7822 : n7862;
  /* TG68K_FPU_ALU.vhd:603:65  */
  assign n7898 = n7808 ? 15'b000000000000001 : n7863;
  /* TG68K_FPU_ALU.vhd:598:65  */
  assign n7899 = n7807 ? sign_a : n7890;
  /* TG68K_FPU_ALU.vhd:598:65  */
  assign n7900 = n7807 ? exp_a : n7891;
  /* TG68K_FPU_ALU.vhd:598:65  */
  assign n7901 = n7807 ? mant_a : n7892;
  /* TG68K_FPU_ALU.vhd:598:65  */
  assign n7902 = n7807 ? mant_sum : n7893;
  /* TG68K_FPU_ALU.vhd:598:65  */
  assign n7904 = n7807 ? mant_a_aligned : n7895;
  /* TG68K_FPU_ALU.vhd:598:65  */
  assign n7905 = n7807 ? mant_b_aligned : n7896;
  /* TG68K_FPU_ALU.vhd:598:65  */
  assign n7906 = n7807 ? exp_larger : n7898;
  /* TG68K_FPU_ALU.vhd:593:65  */
  assign n7907 = n7804 ? n7805 : n7899;
  /* TG68K_FPU_ALU.vhd:593:65  */
  assign n7908 = n7804 ? exp_b : n7900;
  /* TG68K_FPU_ALU.vhd:593:65  */
  assign n7909 = n7804 ? mant_b : n7901;
  /* TG68K_FPU_ALU.vhd:593:65  */
  assign n7910 = n7804 ? mant_sum : n7902;
  /* TG68K_FPU_ALU.vhd:593:65  */
  assign n7912 = n7804 ? mant_a_aligned : n7904;
  /* TG68K_FPU_ALU.vhd:593:65  */
  assign n7913 = n7804 ? mant_b_aligned : n7905;
  /* TG68K_FPU_ALU.vhd:593:65  */
  assign n7914 = n7804 ? exp_larger : n7906;
  /* TG68K_FPU_ALU.vhd:588:65  */
  assign n7915 = is_inf_b ? n7802 : n7907;
  /* TG68K_FPU_ALU.vhd:588:65  */
  assign n7917 = is_inf_b ? 15'b111111111111111 : n7908;
  /* TG68K_FPU_ALU.vhd:588:65  */
  assign n7919 = is_inf_b ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7909;
  /* TG68K_FPU_ALU.vhd:588:65  */
  assign n7920 = is_inf_b ? mant_sum : n7910;
  /* TG68K_FPU_ALU.vhd:588:65  */
  assign n7922 = is_inf_b ? mant_a_aligned : n7912;
  /* TG68K_FPU_ALU.vhd:588:65  */
  assign n7923 = is_inf_b ? mant_b_aligned : n7913;
  /* TG68K_FPU_ALU.vhd:588:65  */
  assign n7924 = is_inf_b ? exp_larger : n7914;
  /* TG68K_FPU_ALU.vhd:583:65  */
  assign n7925 = is_inf_a ? sign_a : n7915;
  /* TG68K_FPU_ALU.vhd:583:65  */
  assign n7927 = is_inf_a ? 15'b111111111111111 : n7917;
  /* TG68K_FPU_ALU.vhd:583:65  */
  assign n7929 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7919;
  /* TG68K_FPU_ALU.vhd:583:65  */
  assign n7930 = is_inf_a ? mant_sum : n7920;
  /* TG68K_FPU_ALU.vhd:583:65  */
  assign n7932 = is_inf_a ? mant_a_aligned : n7922;
  /* TG68K_FPU_ALU.vhd:583:65  */
  assign n7933 = is_inf_a ? mant_b_aligned : n7923;
  /* TG68K_FPU_ALU.vhd:583:65  */
  assign n7934 = is_inf_a ? exp_larger : n7924;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7935 = n7793 ? n7796 : n7925;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7937 = n7793 ? 15'b111111111111111 : n7927;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7938 = n7793 ? n7799 : n7929;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7939 = n7793 ? mant_sum : n7930;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7941 = n7793 ? mant_a_aligned : n7932;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7942 = n7793 ? mant_b_aligned : n7933;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7943 = n7793 ? exp_larger : n7934;
  /* TG68K_FPU_ALU.vhd:569:65  */
  assign n7944 = n7794 & n7793;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7946 = n7792 ? 1'b0 : n7935;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7948 = n7792 ? 15'b111111111111111 : n7937;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7950 = n7792 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n7938;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7951 = n7792 ? mant_sum : n7939;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7953 = n7792 ? mant_a_aligned : n7941;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7954 = n7792 ? mant_b_aligned : n7942;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7955 = n7792 ? exp_larger : n7943;
  /* TG68K_FPU_ALU.vhd:563:65  */
  assign n7957 = n7792 ? 1'b1 : n7801;
  /* TG68K_FPU_ALU.vhd:561:57  */
  assign n7959 = operation_code == 7'b0101000;
  /* TG68K_FPU_ALU.vhd:699:87  */
  assign n7960 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:700:83  */
  assign n7961 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:706:87  */
  assign n7962 = is_zero_b & is_inf_a;
  /* TG68K_FPU_ALU.vhd:706:128  */
  assign n7963 = is_inf_b & is_zero_a;
  /* TG68K_FPU_ALU.vhd:706:108  */
  assign n7964 = n7962 | n7963;
  /* TG68K_FPU_ALU.vhd:712:86  */
  assign n7965 = is_inf_a | is_inf_b;
  /* TG68K_FPU_ALU.vhd:716:87  */
  assign n7966 = is_zero_a | is_zero_b;
  /* TG68K_FPU_ALU.vhd:722:120  */
  assign n7967 = exp_a + exp_b;
  /* TG68K_FPU_ALU.vhd:722:138  */
  assign n7969 = n7967 - 15'b011111111111111;
  /* TG68K_FPU_ALU.vhd:727:135  */
  assign n7970 = {64'b0, mant_a};  //  uext
  /* TG68K_FPU_ALU.vhd:727:135  */
  assign n7971 = {64'b0, mant_b};  //  uext
  /* TG68K_FPU_ALU.vhd:727:135  */
  assign n7972 = n7970 * n7971; // umul
  /* TG68K_FPU_ALU.vhd:729:87  */
  assign n7973 = mult_result[127]; // extract
  /* TG68K_FPU_ALU.vhd:731:133  */
  assign n7975 = exp_result + 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:732:107  */
  assign n7976 = mult_result[126:63]; // extract
  /* TG68K_FPU_ALU.vhd:735:107  */
  assign n7977 = mult_result[125:62]; // extract
  /* TG68K_FPU_ALU.vhd:729:73  */
  assign n7978 = n7973 ? n7975 : n7969;
  /* TG68K_FPU_ALU.vhd:729:73  */
  assign n7979 = n7973 ? n7976 : n7977;
  /* TG68K_FPU_ALU.vhd:738:87  */
  assign n7980 = mult_result[61:0]; // extract
  /* TG68K_FPU_ALU.vhd:738:101  */
  assign n7982 = n7980 != 62'b00000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:738:73  */
  assign n7984 = n7982 ? 1'b1 : flags_inexact;
  /* TG68K_FPU_ALU.vhd:716:65  */
  assign n7986 = n7966 ? 15'b000000000000000 : n7978;
  /* TG68K_FPU_ALU.vhd:716:65  */
  assign n7988 = n7966 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7979;
  /* TG68K_FPU_ALU.vhd:716:65  */
  assign n7989 = n7966 ? mult_result : n7972;
  /* TG68K_FPU_ALU.vhd:716:65  */
  assign n7990 = n7966 ? flags_inexact : n7984;
  /* TG68K_FPU_ALU.vhd:712:65  */
  assign n7992 = n7965 ? 15'b111111111111111 : n7986;
  /* TG68K_FPU_ALU.vhd:712:65  */
  assign n7994 = n7965 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n7988;
  /* TG68K_FPU_ALU.vhd:712:65  */
  assign n7995 = n7965 ? mult_result : n7989;
  /* TG68K_FPU_ALU.vhd:712:65  */
  assign n7996 = n7965 ? flags_inexact : n7990;
  /* TG68K_FPU_ALU.vhd:706:65  */
  assign n7998 = n7964 ? 1'b0 : n7960;
  /* TG68K_FPU_ALU.vhd:706:65  */
  assign n8000 = n7964 ? 15'b111111111111111 : n7992;
  /* TG68K_FPU_ALU.vhd:706:65  */
  assign n8002 = n7964 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n7994;
  /* TG68K_FPU_ALU.vhd:706:65  */
  assign n8003 = n7964 ? mult_result : n7995;
  /* TG68K_FPU_ALU.vhd:706:65  */
  assign n8004 = n7964 ? flags_inexact : n7996;
  /* TG68K_FPU_ALU.vhd:706:65  */
  assign n8006 = n7964 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:700:65  */
  assign n8008 = n7961 ? 1'b0 : n7998;
  /* TG68K_FPU_ALU.vhd:700:65  */
  assign n8010 = n7961 ? 15'b111111111111111 : n8000;
  /* TG68K_FPU_ALU.vhd:700:65  */
  assign n8012 = n7961 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n8002;
  /* TG68K_FPU_ALU.vhd:700:65  */
  assign n8013 = n7961 ? mult_result : n8003;
  /* TG68K_FPU_ALU.vhd:700:65  */
  assign n8014 = n7961 ? flags_inexact : n8004;
  /* TG68K_FPU_ALU.vhd:700:65  */
  assign n8016 = n7961 ? 1'b1 : n8006;
  /* TG68K_FPU_ALU.vhd:697:57  */
  assign n8018 = operation_code == 7'b0100011;
  /* TG68K_FPU_ALU.vhd:746:87  */
  assign n8019 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:747:83  */
  assign n8020 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:753:87  */
  assign n8021 = is_inf_b & is_inf_a;
  /* TG68K_FPU_ALU.vhd:753:127  */
  assign n8022 = is_zero_b & is_zero_a;
  /* TG68K_FPU_ALU.vhd:753:107  */
  assign n8023 = n8021 | n8022;
  /* TG68K_FPU_ALU.vhd:759:91  */
  assign n8024 = ~is_zero_a;
  /* TG68K_FPU_ALU.vhd:759:87  */
  assign n8025 = n8024 & is_zero_b;
  /* TG68K_FPU_ALU.vhd:762:95  */
  assign n8026 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:765:93  */
  assign n8027 = ~is_zero_a;
  /* TG68K_FPU_ALU.vhd:765:89  */
  assign n8028 = n8027 & is_denorm_b;
  /* TG68K_FPU_ALU.vhd:770:95  */
  assign n8033 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:772:82  */
  assign n8034 = mant_b[63:32]; // extract
  /* TG68K_FPU_ALU.vhd:772:97  */
  assign n8036 = n8034 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:779:128  */
  assign n8038 = exp_a - 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:779:149  */
  assign n8040 = n8038 + 15'b011111111111111;
  /* TG68K_FPU_ALU.vhd:780:103  */
  assign n8041 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:772:73  */
  assign n8042 = n8036 ? n8033 : n8041;
  /* TG68K_FPU_ALU.vhd:772:73  */
  assign n8044 = n8036 ? 15'b111111111111111 : n8040;
  /* TG68K_FPU_ALU.vhd:772:73  */
  assign n8046 = n8036 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : mant_result;
  /* TG68K_FPU_ALU.vhd:765:65  */
  assign n8050 = n8095 ? 1'b1 : flags_overflow;
  /* TG68K_FPU_ALU.vhd:797:120  */
  assign n8051 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:797:138  */
  assign n8053 = n8051 + 15'b011111111111111;
  /* TG68K_FPU_ALU.vhd:803:82  */
  assign n8054 = mant_b[63:32]; // extract
  /* TG68K_FPU_ALU.vhd:803:97  */
  assign n8056 = n8054 != 32'b00000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:806:89  */
  assign n8058 = mant_a << 31'b0000000000000000000000000100000;
  /* TG68K_FPU_ALU.vhd:806:139  */
  assign n8059 = mant_b[63:32]; // extract
  /* TG68K_FPU_ALU.vhd:806:122  */
  assign n8060 = {32'b0, n8059};  //  uext
  /* TG68K_FPU_ALU.vhd:806:122  */
  assign n8061 = n8058 / n8060; // udiv
  /* TG68K_FPU_ALU.vhd:808:85  */
  assign n8062 = mant_b[63:16]; // extract
  /* TG68K_FPU_ALU.vhd:808:100  */
  assign n8064 = n8062 != 48'b000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:811:89  */
  assign n8066 = mant_a << 31'b0000000000000000000000000010000;
  /* TG68K_FPU_ALU.vhd:811:139  */
  assign n8067 = mant_b[63:16]; // extract
  /* TG68K_FPU_ALU.vhd:811:122  */
  assign n8068 = {16'b0, n8067};  //  uext
  /* TG68K_FPU_ALU.vhd:811:122  */
  assign n8069 = n8066 / n8068; // udiv
  /* TG68K_FPU_ALU.vhd:816:123  */
  assign n8070 = mant_b[63:1]; // extract
  /* TG68K_FPU_ALU.vhd:816:106  */
  assign n8071 = {1'b0, n8070};  //  uext
  /* TG68K_FPU_ALU.vhd:816:106  */
  assign n8072 = mant_a / n8071; // udiv
  /* TG68K_FPU_ALU.vhd:808:73  */
  assign n8073 = n8064 ? n8069 : n8072;
  /* TG68K_FPU_ALU.vhd:803:73  */
  assign n8074 = n8056 ? n8061 : n8073;
  /* TG68K_FPU_ALU.vhd:791:65  */
  assign n8076 = is_zero_a ? 15'b000000000000000 : n8053;
  /* TG68K_FPU_ALU.vhd:791:65  */
  assign n8078 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n8074;
  /* TG68K_FPU_ALU.vhd:791:65  */
  assign n8080 = is_zero_a ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:787:65  */
  assign n8082 = is_inf_b ? 15'b000000000000000 : n8076;
  /* TG68K_FPU_ALU.vhd:787:65  */
  assign n8084 = is_inf_b ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n8078;
  /* TG68K_FPU_ALU.vhd:787:65  */
  assign n8085 = is_inf_b ? flags_inexact : n8080;
  /* TG68K_FPU_ALU.vhd:783:65  */
  assign n8087 = is_inf_a ? 15'b111111111111111 : n8082;
  /* TG68K_FPU_ALU.vhd:783:65  */
  assign n8089 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n8084;
  /* TG68K_FPU_ALU.vhd:783:65  */
  assign n8090 = is_inf_a ? flags_inexact : n8085;
  /* TG68K_FPU_ALU.vhd:765:65  */
  assign n8091 = n8028 ? n8042 : n8019;
  /* TG68K_FPU_ALU.vhd:765:65  */
  assign n8092 = n8028 ? n8044 : n8087;
  /* TG68K_FPU_ALU.vhd:765:65  */
  assign n8093 = n8028 ? n8046 : n8089;
  /* TG68K_FPU_ALU.vhd:765:65  */
  assign n8095 = n8036 & n8028;
  /* TG68K_FPU_ALU.vhd:765:65  */
  assign n8096 = n8028 ? flags_inexact : n8090;
  /* TG68K_FPU_ALU.vhd:759:65  */
  assign n8097 = n8025 ? n8026 : n8091;
  /* TG68K_FPU_ALU.vhd:759:65  */
  assign n8099 = n8025 ? 15'b111111111111111 : n8092;
  /* TG68K_FPU_ALU.vhd:759:65  */
  assign n8101 = n8025 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n8093;
  /* TG68K_FPU_ALU.vhd:759:65  */
  assign n8103 = n8025 ? flags_overflow : n8050;
  /* TG68K_FPU_ALU.vhd:759:65  */
  assign n8104 = n8025 ? flags_inexact : n8096;
  /* TG68K_FPU_ALU.vhd:759:65  */
  assign n8106 = n8025 ? 1'b1 : flags_div_by_zero;
  /* TG68K_FPU_ALU.vhd:753:65  */
  assign n8108 = n8023 ? 1'b0 : n8097;
  /* TG68K_FPU_ALU.vhd:753:65  */
  assign n8110 = n8023 ? 15'b111111111111111 : n8099;
  /* TG68K_FPU_ALU.vhd:753:65  */
  assign n8112 = n8023 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n8101;
  /* TG68K_FPU_ALU.vhd:753:65  */
  assign n8114 = n8023 ? flags_overflow : n8103;
  /* TG68K_FPU_ALU.vhd:753:65  */
  assign n8115 = n8023 ? flags_inexact : n8104;
  /* TG68K_FPU_ALU.vhd:753:65  */
  assign n8117 = n8023 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:753:65  */
  assign n8118 = n8023 ? flags_div_by_zero : n8106;
  /* TG68K_FPU_ALU.vhd:747:65  */
  assign n8120 = n8020 ? 1'b0 : n8108;
  /* TG68K_FPU_ALU.vhd:747:65  */
  assign n8122 = n8020 ? 15'b111111111111111 : n8110;
  /* TG68K_FPU_ALU.vhd:747:65  */
  assign n8124 = n8020 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n8112;
  /* TG68K_FPU_ALU.vhd:747:65  */
  assign n8126 = n8020 ? flags_overflow : n8114;
  /* TG68K_FPU_ALU.vhd:747:65  */
  assign n8127 = n8020 ? flags_inexact : n8115;
  /* TG68K_FPU_ALU.vhd:747:65  */
  assign n8129 = n8020 ? 1'b1 : n8117;
  /* TG68K_FPU_ALU.vhd:747:65  */
  assign n8130 = n8020 ? flags_div_by_zero : n8118;
  /* TG68K_FPU_ALU.vhd:744:57  */
  assign n8132 = operation_code == 7'b0100000;
  /* TG68K_FPU_ALU.vhd:832:102  */
  assign n8134 = operation_code == 7'b0111000;
  /* TG68K_FPU_ALU.vhd:832:112  */
  assign n8135 = is_nan_b & n8134;
  /* TG68K_FPU_ALU.vhd:832:83  */
  assign n8136 = is_nan_a | n8135;
  /* TG68K_FPU_ALU.vhd:835:107  */
  assign n8138 = operation_code == 7'b0111010;
  /* TG68K_FPU_ALU.vhd:835:117  */
  assign n8139 = n8138 | is_zero_b;
  /* TG68K_FPU_ALU.vhd:835:87  */
  assign n8140 = n8139 & is_zero_a;
  /* TG68K_FPU_ALU.vhd:838:86  */
  assign n8142 = operation_code == 7'b0111010;
  /* TG68K_FPU_ALU.vhd:843:81  */
  assign n8145 = sign_a ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:846:96  */
  assign n8146 = ~is_zero_a;
  /* TG68K_FPU_ALU.vhd:846:92  */
  assign n8147 = n8146 & sign_a;
  /* TG68K_FPU_ALU.vhd:846:73  */
  assign n8150 = n8147 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:840:73  */
  assign n8151 = is_inf_a ? n8145 : n8150;
  /* TG68K_FPU_ALU.vhd:853:83  */
  assign n8152 = sign_a != sign_b;
  /* TG68K_FPU_ALU.vhd:855:81  */
  assign n8155 = sign_a ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:859:85  */
  assign n8156 = exp_a == exp_b;
  /* TG68K_FPU_ALU.vhd:859:104  */
  assign n8157 = mant_a == mant_b;
  /* TG68K_FPU_ALU.vhd:859:93  */
  assign n8158 = n8157 & n8156;
  /* TG68K_FPU_ALU.vhd:861:95  */
  assign n8159 = {exp_a, mant_a};
  /* TG68K_FPU_ALU.vhd:861:122  */
  assign n8160 = {exp_b, mant_b};
  /* TG68K_FPU_ALU.vhd:861:105  */
  assign n8161 = $unsigned(n8159) < $unsigned(n8160);
  /* TG68K_FPU_ALU.vhd:861:133  */
  assign n8162 = n8161 ^ sign_a;
  /* TG68K_FPU_ALU.vhd:861:73  */
  assign n8165 = n8162 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:859:73  */
  assign n8167 = n8158 ? 1'b0 : n8165;
  /* TG68K_FPU_ALU.vhd:853:73  */
  assign n8168 = n8152 ? n8155 : n8167;
  /* TG68K_FPU_ALU.vhd:838:65  */
  assign n8169 = n8142 ? n8151 : n8168;
  /* TG68K_FPU_ALU.vhd:835:65  */
  assign n8171 = n8140 ? 1'b0 : n8169;
  /* TG68K_FPU_ALU.vhd:832:65  */
  assign n8173 = n8136 ? 1'b0 : n8171;
  /* TG68K_FPU_ALU.vhd:832:65  */
  assign n8176 = n8136 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:825:57  */
  assign n8178 = operation_code == 7'b0111000;
  /* TG68K_FPU_ALU.vhd:825:70  */
  assign n8180 = operation_code == 7'b0111010;
  /* TG68K_FPU_ALU.vhd:825:70  */
  assign n8181 = n8178 | n8180;
  /* TG68K_FPU_ALU.vhd:887:77  */
  assign n8183 = $unsigned(exp_a) < $unsigned(15'b011111111111111);
  /* TG68K_FPU_ALU.vhd:889:82  */
  assign n8185 = exp_a == 15'b011111111111110;
  /* TG68K_FPU_ALU.vhd:889:135  */
  assign n8186 = mant_a[63]; // extract
  /* TG68K_FPU_ALU.vhd:889:125  */
  assign n8187 = n8186 & n8185;
  /* TG68K_FPU_ALU.vhd:889:73  */
  assign n8190 = n8187 ? 15'b011111111111111 : 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:889:73  */
  assign n8193 = n8187 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:902:85  */
  assign n8194 = {16'b0, exp_a};  //  uext
  /* TG68K_FPU_ALU.vhd:902:113  */
  assign n8195 = {1'b0, n8194};  //  uext
  /* TG68K_FPU_ALU.vhd:902:113  */
  assign n8197 = n8195 - 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:903:85  */
  assign n8199 = $signed(n8197) >= $signed(32'b00000000000000000000000000111111);
  /* TG68K_FPU_ALU.vhd:913:93  */
  assign n8201 = $signed(n8197) <= $signed(32'b00000000000000000000000000111111);
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8203 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8205 = $signed(32'b00000000000000000000000000000000) < $signed(n8203);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8207 = mant_a[0]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8208 = n8205 ? 1'b0 : n8207;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8210 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8212 = $signed(32'b00000000000000000000000000000001) < $signed(n8210);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8214 = mant_a[1]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8215 = n8212 ? 1'b0 : n8214;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8217 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8219 = $signed(32'b00000000000000000000000000000010) < $signed(n8217);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8221 = mant_a[2]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8222 = n8219 ? 1'b0 : n8221;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8224 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8226 = $signed(32'b00000000000000000000000000000011) < $signed(n8224);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8228 = mant_a[3]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8229 = n8226 ? 1'b0 : n8228;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8231 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8233 = $signed(32'b00000000000000000000000000000100) < $signed(n8231);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8235 = mant_a[4]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8236 = n8233 ? 1'b0 : n8235;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8238 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8240 = $signed(32'b00000000000000000000000000000101) < $signed(n8238);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8242 = mant_a[5]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8243 = n8240 ? 1'b0 : n8242;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8245 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8247 = $signed(32'b00000000000000000000000000000110) < $signed(n8245);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8249 = mant_a[6]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8250 = n8247 ? 1'b0 : n8249;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8252 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8254 = $signed(32'b00000000000000000000000000000111) < $signed(n8252);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8256 = mant_a[7]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8257 = n8254 ? 1'b0 : n8256;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8259 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8261 = $signed(32'b00000000000000000000000000001000) < $signed(n8259);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8263 = mant_a[8]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8264 = n8261 ? 1'b0 : n8263;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8266 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8268 = $signed(32'b00000000000000000000000000001001) < $signed(n8266);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8270 = mant_a[9]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8271 = n8268 ? 1'b0 : n8270;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8273 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8275 = $signed(32'b00000000000000000000000000001010) < $signed(n8273);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8277 = mant_a[10]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8278 = n8275 ? 1'b0 : n8277;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8280 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8282 = $signed(32'b00000000000000000000000000001011) < $signed(n8280);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8284 = mant_a[11]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8285 = n8282 ? 1'b0 : n8284;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8287 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8289 = $signed(32'b00000000000000000000000000001100) < $signed(n8287);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8291 = mant_a[12]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8292 = n8289 ? 1'b0 : n8291;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8294 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8296 = $signed(32'b00000000000000000000000000001101) < $signed(n8294);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8298 = mant_a[13]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8299 = n8296 ? 1'b0 : n8298;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8301 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8303 = $signed(32'b00000000000000000000000000001110) < $signed(n8301);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8305 = mant_a[14]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8306 = n8303 ? 1'b0 : n8305;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8308 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8310 = $signed(32'b00000000000000000000000000001111) < $signed(n8308);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8312 = mant_a[15]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8313 = n8310 ? 1'b0 : n8312;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8315 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8317 = $signed(32'b00000000000000000000000000010000) < $signed(n8315);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8319 = mant_a[16]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8320 = n8317 ? 1'b0 : n8319;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8322 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8324 = $signed(32'b00000000000000000000000000010001) < $signed(n8322);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8326 = mant_a[17]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8327 = n8324 ? 1'b0 : n8326;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8329 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8331 = $signed(32'b00000000000000000000000000010010) < $signed(n8329);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8333 = mant_a[18]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8334 = n8331 ? 1'b0 : n8333;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8336 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8338 = $signed(32'b00000000000000000000000000010011) < $signed(n8336);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8340 = mant_a[19]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8341 = n8338 ? 1'b0 : n8340;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8343 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8345 = $signed(32'b00000000000000000000000000010100) < $signed(n8343);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8347 = mant_a[20]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8348 = n8345 ? 1'b0 : n8347;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8350 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8352 = $signed(32'b00000000000000000000000000010101) < $signed(n8350);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8354 = mant_a[21]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8355 = n8352 ? 1'b0 : n8354;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8357 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8359 = $signed(32'b00000000000000000000000000010110) < $signed(n8357);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8361 = mant_a[22]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8362 = n8359 ? 1'b0 : n8361;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8364 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8366 = $signed(32'b00000000000000000000000000010111) < $signed(n8364);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8368 = mant_a[23]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8369 = n8366 ? 1'b0 : n8368;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8371 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8373 = $signed(32'b00000000000000000000000000011000) < $signed(n8371);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8375 = mant_a[24]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8376 = n8373 ? 1'b0 : n8375;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8378 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8380 = $signed(32'b00000000000000000000000000011001) < $signed(n8378);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8382 = mant_a[25]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8383 = n8380 ? 1'b0 : n8382;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8385 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8387 = $signed(32'b00000000000000000000000000011010) < $signed(n8385);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8389 = mant_a[26]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8390 = n8387 ? 1'b0 : n8389;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8392 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8394 = $signed(32'b00000000000000000000000000011011) < $signed(n8392);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8396 = mant_a[27]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8397 = n8394 ? 1'b0 : n8396;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8399 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8401 = $signed(32'b00000000000000000000000000011100) < $signed(n8399);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8403 = mant_a[28]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8404 = n8401 ? 1'b0 : n8403;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8406 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8408 = $signed(32'b00000000000000000000000000011101) < $signed(n8406);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8410 = mant_a[29]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8411 = n8408 ? 1'b0 : n8410;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8413 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8415 = $signed(32'b00000000000000000000000000011110) < $signed(n8413);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8417 = mant_a[30]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8418 = n8415 ? 1'b0 : n8417;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8420 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8422 = $signed(32'b00000000000000000000000000011111) < $signed(n8420);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8424 = mant_a[31]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8425 = n8422 ? 1'b0 : n8424;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8427 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8429 = $signed(32'b00000000000000000000000000100000) < $signed(n8427);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8431 = mant_a[32]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8432 = n8429 ? 1'b0 : n8431;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8434 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8436 = $signed(32'b00000000000000000000000000100001) < $signed(n8434);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8438 = mant_a[33]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8439 = n8436 ? 1'b0 : n8438;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8441 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8443 = $signed(32'b00000000000000000000000000100010) < $signed(n8441);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8445 = mant_a[34]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8446 = n8443 ? 1'b0 : n8445;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8448 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8450 = $signed(32'b00000000000000000000000000100011) < $signed(n8448);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8452 = mant_a[35]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8453 = n8450 ? 1'b0 : n8452;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8455 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8457 = $signed(32'b00000000000000000000000000100100) < $signed(n8455);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8459 = mant_a[36]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8460 = n8457 ? 1'b0 : n8459;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8462 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8464 = $signed(32'b00000000000000000000000000100101) < $signed(n8462);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8466 = mant_a[37]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8467 = n8464 ? 1'b0 : n8466;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8469 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8471 = $signed(32'b00000000000000000000000000100110) < $signed(n8469);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8473 = mant_a[38]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8474 = n8471 ? 1'b0 : n8473;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8476 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8478 = $signed(32'b00000000000000000000000000100111) < $signed(n8476);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8480 = mant_a[39]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8481 = n8478 ? 1'b0 : n8480;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8483 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8485 = $signed(32'b00000000000000000000000000101000) < $signed(n8483);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8487 = mant_a[40]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8488 = n8485 ? 1'b0 : n8487;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8490 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8492 = $signed(32'b00000000000000000000000000101001) < $signed(n8490);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8494 = mant_a[41]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8495 = n8492 ? 1'b0 : n8494;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8497 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8499 = $signed(32'b00000000000000000000000000101010) < $signed(n8497);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8501 = mant_a[42]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8502 = n8499 ? 1'b0 : n8501;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8504 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8506 = $signed(32'b00000000000000000000000000101011) < $signed(n8504);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8508 = mant_a[43]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8509 = n8506 ? 1'b0 : n8508;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8511 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8513 = $signed(32'b00000000000000000000000000101100) < $signed(n8511);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8515 = mant_a[44]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8516 = n8513 ? 1'b0 : n8515;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8518 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8520 = $signed(32'b00000000000000000000000000101101) < $signed(n8518);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8522 = mant_a[45]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8523 = n8520 ? 1'b0 : n8522;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8525 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8527 = $signed(32'b00000000000000000000000000101110) < $signed(n8525);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8529 = mant_a[46]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8530 = n8527 ? 1'b0 : n8529;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8532 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8534 = $signed(32'b00000000000000000000000000101111) < $signed(n8532);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8536 = mant_a[47]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8537 = n8534 ? 1'b0 : n8536;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8539 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8541 = $signed(32'b00000000000000000000000000110000) < $signed(n8539);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8543 = mant_a[48]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8544 = n8541 ? 1'b0 : n8543;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8546 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8548 = $signed(32'b00000000000000000000000000110001) < $signed(n8546);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8550 = mant_a[49]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8551 = n8548 ? 1'b0 : n8550;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8553 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8555 = $signed(32'b00000000000000000000000000110010) < $signed(n8553);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8557 = mant_a[50]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8558 = n8555 ? 1'b0 : n8557;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8560 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8562 = $signed(32'b00000000000000000000000000110011) < $signed(n8560);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8564 = mant_a[51]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8565 = n8562 ? 1'b0 : n8564;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8567 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8569 = $signed(32'b00000000000000000000000000110100) < $signed(n8567);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8571 = mant_a[52]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8572 = n8569 ? 1'b0 : n8571;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8574 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8576 = $signed(32'b00000000000000000000000000110101) < $signed(n8574);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8578 = mant_a[53]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8579 = n8576 ? 1'b0 : n8578;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8581 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8583 = $signed(32'b00000000000000000000000000110110) < $signed(n8581);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8585 = mant_a[54]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8586 = n8583 ? 1'b0 : n8585;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8588 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8590 = $signed(32'b00000000000000000000000000110111) < $signed(n8588);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8592 = mant_a[55]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8593 = n8590 ? 1'b0 : n8592;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8595 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8597 = $signed(32'b00000000000000000000000000111000) < $signed(n8595);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8599 = mant_a[56]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8600 = n8597 ? 1'b0 : n8599;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8602 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8604 = $signed(32'b00000000000000000000000000111001) < $signed(n8602);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8606 = mant_a[57]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8607 = n8604 ? 1'b0 : n8606;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8609 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8611 = $signed(32'b00000000000000000000000000111010) < $signed(n8609);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8613 = mant_a[58]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8614 = n8611 ? 1'b0 : n8613;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8616 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8618 = $signed(32'b00000000000000000000000000111011) < $signed(n8616);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8620 = mant_a[59]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8621 = n8618 ? 1'b0 : n8620;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8623 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8625 = $signed(32'b00000000000000000000000000111100) < $signed(n8623);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8627 = mant_a[60]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8628 = n8625 ? 1'b0 : n8627;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8630 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8632 = $signed(32'b00000000000000000000000000111101) < $signed(n8630);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8634 = mant_a[61]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8635 = n8632 ? 1'b0 : n8634;
  /* TG68K_FPU_ALU.vhd:915:108  */
  assign n8637 = 32'b00000000000000000000000000111111 - n8197;
  /* TG68K_FPU_ALU.vhd:915:102  */
  assign n8639 = $signed(32'b00000000000000000000000000111110) < $signed(n8637);
  /* TG68K_FPU_ALU.vhd:918:129  */
  assign n8641 = mant_a[62]; // extract
  /* TG68K_FPU_ALU.vhd:915:97  */
  assign n8642 = n8639 ? 1'b0 : n8641;
  /* TG68K_FPU_ALU.vhd:921:114  */
  assign n8643 = mant_a[63]; // extract
  assign n8644 = {n8643, n8642, n8635, n8628, n8621, n8614, n8607, n8600, n8593, n8586, n8579, n8572, n8565, n8558, n8551, n8544, n8537, n8530, n8523, n8516, n8509, n8502, n8495, n8488, n8481, n8474, n8467, n8460, n8453, n8446, n8439, n8432, n8425, n8418, n8411, n8404, n8397, n8390, n8383, n8376, n8369, n8362, n8355, n8348, n8341, n8334, n8327, n8320, n8313, n8306, n8299, n8292, n8285, n8278, n8271, n8264, n8257, n8250, n8243, n8236, n8229, n8222, n8215, n8208};
  /* TG68K_FPU_ALU.vhd:913:81  */
  assign n8645 = n8201 ? n8644 : mant_a;
  /* TG68K_FPU_ALU.vhd:903:73  */
  assign n8646 = n8199 ? mant_a : n8645;
  /* TG68K_FPU_ALU.vhd:887:65  */
  assign n8647 = n8183 ? n8190 : exp_a;
  /* TG68K_FPU_ALU.vhd:887:65  */
  assign n8648 = n8183 ? n8193 : n8646;
  /* TG68K_FPU_ALU.vhd:887:65  */
  assign n8650 = n8183 ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:882:65  */
  assign n8653 = is_zero_a ? 15'b000000000000000 : n8647;
  /* TG68K_FPU_ALU.vhd:882:65  */
  assign n8655 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n8648;
  /* TG68K_FPU_ALU.vhd:882:65  */
  assign n8656 = is_zero_a ? flags_inexact : n8650;
  /* TG68K_FPU_ALU.vhd:877:65  */
  assign n8659 = is_inf_a ? 15'b111111111111111 : n8653;
  /* TG68K_FPU_ALU.vhd:877:65  */
  assign n8661 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n8655;
  /* TG68K_FPU_ALU.vhd:877:65  */
  assign n8662 = is_inf_a ? flags_inexact : n8656;
  /* TG68K_FPU_ALU.vhd:871:65  */
  assign n8665 = is_nan_a ? 1'b0 : sign_a;
  /* TG68K_FPU_ALU.vhd:871:65  */
  assign n8667 = is_nan_a ? 15'b111111111111111 : n8659;
  /* TG68K_FPU_ALU.vhd:871:65  */
  assign n8669 = is_nan_a ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n8661;
  /* TG68K_FPU_ALU.vhd:871:65  */
  assign n8670 = is_nan_a ? flags_inexact : n8662;
  /* TG68K_FPU_ALU.vhd:871:65  */
  assign n8672 = is_nan_a ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:869:57  */
  assign n8675 = operation_code == 7'b0000001;
  /* TG68K_FPU_ALU.vhd:948:77  */
  assign n8677 = $unsigned(exp_a) < $unsigned(15'b011111111111111);
  /* TG68K_FPU_ALU.vhd:955:85  */
  assign n8678 = {16'b0, exp_a};  //  uext
  /* TG68K_FPU_ALU.vhd:955:113  */
  assign n8679 = {1'b0, n8678};  //  uext
  /* TG68K_FPU_ALU.vhd:955:113  */
  assign n8681 = n8679 - 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:956:85  */
  assign n8683 = $signed(n8681) >= $signed(32'b00000000000000000000000000111111);
  /* TG68K_FPU_ALU.vhd:966:93  */
  assign n8685 = $signed(n8681) <= $signed(32'b00000000000000000000000000111111);
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8687 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8689 = $signed(32'b00000000000000000000000000000000) < $signed(n8687);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8691 = mant_a[0]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8692 = n8689 ? 1'b0 : n8691;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8694 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8696 = $signed(32'b00000000000000000000000000000001) < $signed(n8694);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8698 = mant_a[1]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8699 = n8696 ? 1'b0 : n8698;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8701 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8703 = $signed(32'b00000000000000000000000000000010) < $signed(n8701);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8705 = mant_a[2]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8706 = n8703 ? 1'b0 : n8705;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8708 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8710 = $signed(32'b00000000000000000000000000000011) < $signed(n8708);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8712 = mant_a[3]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8713 = n8710 ? 1'b0 : n8712;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8715 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8717 = $signed(32'b00000000000000000000000000000100) < $signed(n8715);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8719 = mant_a[4]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8720 = n8717 ? 1'b0 : n8719;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8722 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8724 = $signed(32'b00000000000000000000000000000101) < $signed(n8722);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8726 = mant_a[5]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8727 = n8724 ? 1'b0 : n8726;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8729 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8731 = $signed(32'b00000000000000000000000000000110) < $signed(n8729);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8733 = mant_a[6]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8734 = n8731 ? 1'b0 : n8733;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8736 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8738 = $signed(32'b00000000000000000000000000000111) < $signed(n8736);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8740 = mant_a[7]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8741 = n8738 ? 1'b0 : n8740;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8743 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8745 = $signed(32'b00000000000000000000000000001000) < $signed(n8743);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8747 = mant_a[8]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8748 = n8745 ? 1'b0 : n8747;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8750 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8752 = $signed(32'b00000000000000000000000000001001) < $signed(n8750);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8754 = mant_a[9]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8755 = n8752 ? 1'b0 : n8754;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8757 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8759 = $signed(32'b00000000000000000000000000001010) < $signed(n8757);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8761 = mant_a[10]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8762 = n8759 ? 1'b0 : n8761;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8764 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8766 = $signed(32'b00000000000000000000000000001011) < $signed(n8764);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8768 = mant_a[11]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8769 = n8766 ? 1'b0 : n8768;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8771 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8773 = $signed(32'b00000000000000000000000000001100) < $signed(n8771);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8775 = mant_a[12]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8776 = n8773 ? 1'b0 : n8775;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8778 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8780 = $signed(32'b00000000000000000000000000001101) < $signed(n8778);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8782 = mant_a[13]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8783 = n8780 ? 1'b0 : n8782;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8785 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8787 = $signed(32'b00000000000000000000000000001110) < $signed(n8785);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8789 = mant_a[14]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8790 = n8787 ? 1'b0 : n8789;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8792 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8794 = $signed(32'b00000000000000000000000000001111) < $signed(n8792);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8796 = mant_a[15]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8797 = n8794 ? 1'b0 : n8796;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8799 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8801 = $signed(32'b00000000000000000000000000010000) < $signed(n8799);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8803 = mant_a[16]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8804 = n8801 ? 1'b0 : n8803;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8806 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8808 = $signed(32'b00000000000000000000000000010001) < $signed(n8806);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8810 = mant_a[17]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8811 = n8808 ? 1'b0 : n8810;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8813 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8815 = $signed(32'b00000000000000000000000000010010) < $signed(n8813);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8817 = mant_a[18]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8818 = n8815 ? 1'b0 : n8817;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8820 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8822 = $signed(32'b00000000000000000000000000010011) < $signed(n8820);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8824 = mant_a[19]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8825 = n8822 ? 1'b0 : n8824;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8827 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8829 = $signed(32'b00000000000000000000000000010100) < $signed(n8827);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8831 = mant_a[20]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8832 = n8829 ? 1'b0 : n8831;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8834 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8836 = $signed(32'b00000000000000000000000000010101) < $signed(n8834);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8838 = mant_a[21]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8839 = n8836 ? 1'b0 : n8838;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8841 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8843 = $signed(32'b00000000000000000000000000010110) < $signed(n8841);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8845 = mant_a[22]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8846 = n8843 ? 1'b0 : n8845;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8848 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8850 = $signed(32'b00000000000000000000000000010111) < $signed(n8848);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8852 = mant_a[23]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8853 = n8850 ? 1'b0 : n8852;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8855 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8857 = $signed(32'b00000000000000000000000000011000) < $signed(n8855);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8859 = mant_a[24]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8860 = n8857 ? 1'b0 : n8859;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8862 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8864 = $signed(32'b00000000000000000000000000011001) < $signed(n8862);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8866 = mant_a[25]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8867 = n8864 ? 1'b0 : n8866;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8869 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8871 = $signed(32'b00000000000000000000000000011010) < $signed(n8869);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8873 = mant_a[26]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8874 = n8871 ? 1'b0 : n8873;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8876 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8878 = $signed(32'b00000000000000000000000000011011) < $signed(n8876);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8880 = mant_a[27]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8881 = n8878 ? 1'b0 : n8880;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8883 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8885 = $signed(32'b00000000000000000000000000011100) < $signed(n8883);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8887 = mant_a[28]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8888 = n8885 ? 1'b0 : n8887;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8890 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8892 = $signed(32'b00000000000000000000000000011101) < $signed(n8890);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8894 = mant_a[29]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8895 = n8892 ? 1'b0 : n8894;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8897 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8899 = $signed(32'b00000000000000000000000000011110) < $signed(n8897);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8901 = mant_a[30]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8902 = n8899 ? 1'b0 : n8901;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8904 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8906 = $signed(32'b00000000000000000000000000011111) < $signed(n8904);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8908 = mant_a[31]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8909 = n8906 ? 1'b0 : n8908;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8911 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8913 = $signed(32'b00000000000000000000000000100000) < $signed(n8911);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8915 = mant_a[32]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8916 = n8913 ? 1'b0 : n8915;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8918 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8920 = $signed(32'b00000000000000000000000000100001) < $signed(n8918);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8922 = mant_a[33]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8923 = n8920 ? 1'b0 : n8922;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8925 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8927 = $signed(32'b00000000000000000000000000100010) < $signed(n8925);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8929 = mant_a[34]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8930 = n8927 ? 1'b0 : n8929;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8932 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8934 = $signed(32'b00000000000000000000000000100011) < $signed(n8932);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8936 = mant_a[35]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8937 = n8934 ? 1'b0 : n8936;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8939 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8941 = $signed(32'b00000000000000000000000000100100) < $signed(n8939);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8943 = mant_a[36]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8944 = n8941 ? 1'b0 : n8943;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8946 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8948 = $signed(32'b00000000000000000000000000100101) < $signed(n8946);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8950 = mant_a[37]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8951 = n8948 ? 1'b0 : n8950;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8953 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8955 = $signed(32'b00000000000000000000000000100110) < $signed(n8953);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8957 = mant_a[38]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8958 = n8955 ? 1'b0 : n8957;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8960 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8962 = $signed(32'b00000000000000000000000000100111) < $signed(n8960);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8964 = mant_a[39]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8965 = n8962 ? 1'b0 : n8964;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8967 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8969 = $signed(32'b00000000000000000000000000101000) < $signed(n8967);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8971 = mant_a[40]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8972 = n8969 ? 1'b0 : n8971;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8974 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8976 = $signed(32'b00000000000000000000000000101001) < $signed(n8974);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8978 = mant_a[41]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8979 = n8976 ? 1'b0 : n8978;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8981 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8983 = $signed(32'b00000000000000000000000000101010) < $signed(n8981);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8985 = mant_a[42]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8986 = n8983 ? 1'b0 : n8985;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8988 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8990 = $signed(32'b00000000000000000000000000101011) < $signed(n8988);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8992 = mant_a[43]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n8993 = n8990 ? 1'b0 : n8992;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n8995 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n8997 = $signed(32'b00000000000000000000000000101100) < $signed(n8995);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n8999 = mant_a[44]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9000 = n8997 ? 1'b0 : n8999;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9002 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9004 = $signed(32'b00000000000000000000000000101101) < $signed(n9002);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9006 = mant_a[45]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9007 = n9004 ? 1'b0 : n9006;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9009 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9011 = $signed(32'b00000000000000000000000000101110) < $signed(n9009);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9013 = mant_a[46]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9014 = n9011 ? 1'b0 : n9013;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9016 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9018 = $signed(32'b00000000000000000000000000101111) < $signed(n9016);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9020 = mant_a[47]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9021 = n9018 ? 1'b0 : n9020;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9023 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9025 = $signed(32'b00000000000000000000000000110000) < $signed(n9023);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9027 = mant_a[48]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9028 = n9025 ? 1'b0 : n9027;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9030 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9032 = $signed(32'b00000000000000000000000000110001) < $signed(n9030);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9034 = mant_a[49]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9035 = n9032 ? 1'b0 : n9034;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9037 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9039 = $signed(32'b00000000000000000000000000110010) < $signed(n9037);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9041 = mant_a[50]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9042 = n9039 ? 1'b0 : n9041;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9044 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9046 = $signed(32'b00000000000000000000000000110011) < $signed(n9044);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9048 = mant_a[51]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9049 = n9046 ? 1'b0 : n9048;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9051 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9053 = $signed(32'b00000000000000000000000000110100) < $signed(n9051);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9055 = mant_a[52]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9056 = n9053 ? 1'b0 : n9055;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9058 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9060 = $signed(32'b00000000000000000000000000110101) < $signed(n9058);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9062 = mant_a[53]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9063 = n9060 ? 1'b0 : n9062;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9065 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9067 = $signed(32'b00000000000000000000000000110110) < $signed(n9065);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9069 = mant_a[54]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9070 = n9067 ? 1'b0 : n9069;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9072 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9074 = $signed(32'b00000000000000000000000000110111) < $signed(n9072);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9076 = mant_a[55]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9077 = n9074 ? 1'b0 : n9076;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9079 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9081 = $signed(32'b00000000000000000000000000111000) < $signed(n9079);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9083 = mant_a[56]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9084 = n9081 ? 1'b0 : n9083;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9086 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9088 = $signed(32'b00000000000000000000000000111001) < $signed(n9086);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9090 = mant_a[57]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9091 = n9088 ? 1'b0 : n9090;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9093 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9095 = $signed(32'b00000000000000000000000000111010) < $signed(n9093);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9097 = mant_a[58]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9098 = n9095 ? 1'b0 : n9097;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9100 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9102 = $signed(32'b00000000000000000000000000111011) < $signed(n9100);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9104 = mant_a[59]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9105 = n9102 ? 1'b0 : n9104;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9107 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9109 = $signed(32'b00000000000000000000000000111100) < $signed(n9107);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9111 = mant_a[60]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9112 = n9109 ? 1'b0 : n9111;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9114 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9116 = $signed(32'b00000000000000000000000000111101) < $signed(n9114);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9118 = mant_a[61]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9119 = n9116 ? 1'b0 : n9118;
  /* TG68K_FPU_ALU.vhd:968:108  */
  assign n9121 = 32'b00000000000000000000000000111111 - n8681;
  /* TG68K_FPU_ALU.vhd:968:102  */
  assign n9123 = $signed(32'b00000000000000000000000000111110) < $signed(n9121);
  /* TG68K_FPU_ALU.vhd:971:129  */
  assign n9125 = mant_a[62]; // extract
  /* TG68K_FPU_ALU.vhd:968:97  */
  assign n9126 = n9123 ? 1'b0 : n9125;
  /* TG68K_FPU_ALU.vhd:974:114  */
  assign n9127 = mant_a[63]; // extract
  assign n9128 = {n9127, n9126, n9119, n9112, n9105, n9098, n9091, n9084, n9077, n9070, n9063, n9056, n9049, n9042, n9035, n9028, n9021, n9014, n9007, n9000, n8993, n8986, n8979, n8972, n8965, n8958, n8951, n8944, n8937, n8930, n8923, n8916, n8909, n8902, n8895, n8888, n8881, n8874, n8867, n8860, n8853, n8846, n8839, n8832, n8825, n8818, n8811, n8804, n8797, n8790, n8783, n8776, n8769, n8762, n8755, n8748, n8741, n8734, n8727, n8720, n8713, n8706, n8699, n8692};
  /* TG68K_FPU_ALU.vhd:966:81  */
  assign n9129 = n8685 ? n9128 : mant_a;
  /* TG68K_FPU_ALU.vhd:956:73  */
  assign n9130 = n8683 ? mant_a : n9129;
  /* TG68K_FPU_ALU.vhd:948:65  */
  assign n9132 = n8677 ? 15'b000000000000000 : exp_a;
  /* TG68K_FPU_ALU.vhd:948:65  */
  assign n9134 = n8677 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9130;
  /* TG68K_FPU_ALU.vhd:948:65  */
  assign n9136 = n8677 ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:943:65  */
  assign n9139 = is_zero_a ? 15'b000000000000000 : n9132;
  /* TG68K_FPU_ALU.vhd:943:65  */
  assign n9141 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9134;
  /* TG68K_FPU_ALU.vhd:943:65  */
  assign n9142 = is_zero_a ? flags_inexact : n9136;
  /* TG68K_FPU_ALU.vhd:938:65  */
  assign n9145 = is_inf_a ? 15'b111111111111111 : n9139;
  /* TG68K_FPU_ALU.vhd:938:65  */
  assign n9147 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9141;
  /* TG68K_FPU_ALU.vhd:938:65  */
  assign n9148 = is_inf_a ? flags_inexact : n9142;
  /* TG68K_FPU_ALU.vhd:932:65  */
  assign n9151 = is_nan_a ? 1'b0 : sign_a;
  /* TG68K_FPU_ALU.vhd:932:65  */
  assign n9153 = is_nan_a ? 15'b111111111111111 : n9145;
  /* TG68K_FPU_ALU.vhd:932:65  */
  assign n9155 = is_nan_a ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9147;
  /* TG68K_FPU_ALU.vhd:932:65  */
  assign n9156 = is_nan_a ? flags_inexact : n9148;
  /* TG68K_FPU_ALU.vhd:932:65  */
  assign n9158 = is_nan_a ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:930:57  */
  assign n9161 = operation_code == 7'b0000011;
  /* TG68K_FPU_ALU.vhd:985:87  */
  assign n9162 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:986:83  */
  assign n9163 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:992:87  */
  assign n9164 = is_inf_b & is_inf_a;
  /* TG68K_FPU_ALU.vhd:992:127  */
  assign n9165 = is_zero_b & is_zero_a;
  /* TG68K_FPU_ALU.vhd:992:107  */
  assign n9166 = n9164 | n9165;
  /* TG68K_FPU_ALU.vhd:998:91  */
  assign n9167 = ~is_zero_a;
  /* TG68K_FPU_ALU.vhd:998:87  */
  assign n9168 = n9167 & is_zero_b;
  /* TG68K_FPU_ALU.vhd:1017:120  */
  assign n9169 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:1017:138  */
  assign n9171 = n9169 + 15'b011111111111111;
  /* TG68K_FPU_ALU.vhd:1019:83  */
  assign n9172 = mant_a == mant_b;
  /* TG68K_FPU_ALU.vhd:1021:96  */
  assign n9173 = $unsigned(mant_a) > $unsigned(mant_b);
  /* TG68K_FPU_ALU.vhd:1022:90  */
  assign n9174 = mant_b[63:48]; // extract
  /* TG68K_FPU_ALU.vhd:1022:105  */
  assign n9176 = n9174 != 16'b0000000000000000;
  /* TG68K_FPU_ALU.vhd:1024:112  */
  assign n9177 = mant_a[63:32]; // extract
  /* TG68K_FPU_ALU.vhd:1024:128  */
  assign n9178 = {32'b0, n9177};  //  uext
  /* TG68K_FPU_ALU.vhd:1024:128  */
  assign n9180 = $signed(n9178) * $signed(64'b0000000000000000000000000000000000000000000000000000100000000000); // smul
  /* TG68K_FPU_ALU.vhd:1024:152  */
  assign n9181 = mant_b[63:48]; // extract
  /* TG68K_FPU_ALU.vhd:1024:135  */
  assign n9182 = {48'b0, n9181};  //  uext
  /* TG68K_FPU_ALU.vhd:1024:135  */
  assign n9183 = n9180 / n9182; // udiv
  /* TG68K_FPU_ALU.vhd:1022:81  */
  assign n9185 = n9176 ? n9183 : 64'b1111111111111111111111111111111111111111111111111111111111111111;
  /* TG68K_FPU_ALU.vhd:1022:81  */
  assign n9187 = n9176 ? flags_overflow : 1'b1;
  /* TG68K_FPU_ALU.vhd:1031:133  */
  assign n9189 = exp_result - 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:1032:90  */
  assign n9190 = mant_b[63:48]; // extract
  /* TG68K_FPU_ALU.vhd:1032:105  */
  assign n9192 = n9190 != 16'b0000000000000000;
  /* TG68K_FPU_ALU.vhd:1035:112  */
  assign n9193 = mant_a[63:32]; // extract
  /* TG68K_FPU_ALU.vhd:1035:128  */
  assign n9194 = {32'b0, n9193};  //  uext
  /* TG68K_FPU_ALU.vhd:1035:128  */
  assign n9196 = $signed(n9194) * $signed(64'b0000000000000000000000000000000000000000000000000001000000000000); // smul
  /* TG68K_FPU_ALU.vhd:1035:152  */
  assign n9197 = mant_b[63:48]; // extract
  /* TG68K_FPU_ALU.vhd:1035:135  */
  assign n9198 = {48'b0, n9197};  //  uext
  /* TG68K_FPU_ALU.vhd:1035:135  */
  assign n9199 = n9196 / n9198; // udiv
  /* TG68K_FPU_ALU.vhd:1038:110  */
  assign n9200 = mant_a[62:0]; // extract
  /* TG68K_FPU_ALU.vhd:1038:124  */
  assign n9202 = {n9200, 1'b0};
  /* TG68K_FPU_ALU.vhd:1032:81  */
  assign n9203 = n9192 ? n9199 : n9202;
  /* TG68K_FPU_ALU.vhd:1021:73  */
  assign n9204 = n9173 ? n9171 : n9189;
  /* TG68K_FPU_ALU.vhd:1021:73  */
  assign n9205 = n9173 ? n9185 : n9203;
  /* TG68K_FPU_ALU.vhd:1021:73  */
  assign n9206 = n9173 ? n9187 : flags_overflow;
  /* TG68K_FPU_ALU.vhd:1019:73  */
  assign n9207 = n9172 ? n9171 : n9204;
  /* TG68K_FPU_ALU.vhd:1019:73  */
  assign n9209 = n9172 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9205;
  /* TG68K_FPU_ALU.vhd:1019:73  */
  assign n9210 = n9172 ? flags_overflow : n9206;
  assign n9212 = n9209[63:40]; // extract
  /* TG68K_FPU_ALU.vhd:1011:65  */
  assign n9214 = is_zero_a ? 15'b000000000000000 : n9207;
  assign n9215 = {n9212, 40'b0000000000000000000000000000000000000000};
  /* TG68K_FPU_ALU.vhd:1011:65  */
  assign n9217 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9215;
  /* TG68K_FPU_ALU.vhd:1011:65  */
  assign n9218 = is_zero_a ? flags_overflow : n9210;
  /* TG68K_FPU_ALU.vhd:1011:65  */
  assign n9220 = is_zero_a ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:1007:65  */
  assign n9222 = is_inf_b ? 15'b000000000000000 : n9214;
  /* TG68K_FPU_ALU.vhd:1007:65  */
  assign n9224 = is_inf_b ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9217;
  /* TG68K_FPU_ALU.vhd:1007:65  */
  assign n9225 = is_inf_b ? flags_overflow : n9218;
  /* TG68K_FPU_ALU.vhd:1007:65  */
  assign n9226 = is_inf_b ? flags_inexact : n9220;
  /* TG68K_FPU_ALU.vhd:1003:65  */
  assign n9228 = is_inf_a ? 15'b111111111111111 : n9222;
  /* TG68K_FPU_ALU.vhd:1003:65  */
  assign n9230 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9224;
  /* TG68K_FPU_ALU.vhd:1003:65  */
  assign n9231 = is_inf_a ? flags_overflow : n9225;
  /* TG68K_FPU_ALU.vhd:1003:65  */
  assign n9232 = is_inf_a ? flags_inexact : n9226;
  /* TG68K_FPU_ALU.vhd:998:65  */
  assign n9234 = n9168 ? 15'b111111111111111 : n9228;
  /* TG68K_FPU_ALU.vhd:998:65  */
  assign n9236 = n9168 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9230;
  /* TG68K_FPU_ALU.vhd:998:65  */
  assign n9237 = n9168 ? flags_overflow : n9231;
  /* TG68K_FPU_ALU.vhd:998:65  */
  assign n9238 = n9168 ? flags_inexact : n9232;
  /* TG68K_FPU_ALU.vhd:998:65  */
  assign n9240 = n9168 ? 1'b1 : flags_div_by_zero;
  /* TG68K_FPU_ALU.vhd:992:65  */
  assign n9242 = n9166 ? 1'b0 : n9162;
  /* TG68K_FPU_ALU.vhd:992:65  */
  assign n9244 = n9166 ? 15'b111111111111111 : n9234;
  /* TG68K_FPU_ALU.vhd:992:65  */
  assign n9246 = n9166 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9236;
  /* TG68K_FPU_ALU.vhd:992:65  */
  assign n9247 = n9166 ? flags_overflow : n9237;
  /* TG68K_FPU_ALU.vhd:992:65  */
  assign n9248 = n9166 ? flags_inexact : n9238;
  /* TG68K_FPU_ALU.vhd:992:65  */
  assign n9250 = n9166 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:992:65  */
  assign n9251 = n9166 ? flags_div_by_zero : n9240;
  /* TG68K_FPU_ALU.vhd:986:65  */
  assign n9253 = n9163 ? 1'b0 : n9242;
  /* TG68K_FPU_ALU.vhd:986:65  */
  assign n9255 = n9163 ? 15'b111111111111111 : n9244;
  /* TG68K_FPU_ALU.vhd:986:65  */
  assign n9257 = n9163 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9246;
  /* TG68K_FPU_ALU.vhd:986:65  */
  assign n9258 = n9163 ? flags_overflow : n9247;
  /* TG68K_FPU_ALU.vhd:986:65  */
  assign n9259 = n9163 ? flags_inexact : n9248;
  /* TG68K_FPU_ALU.vhd:986:65  */
  assign n9261 = n9163 ? 1'b1 : n9250;
  /* TG68K_FPU_ALU.vhd:986:65  */
  assign n9262 = n9163 ? flags_div_by_zero : n9251;
  /* TG68K_FPU_ALU.vhd:983:57  */
  assign n9264 = operation_code == 7'b0100100;
  /* TG68K_FPU_ALU.vhd:1049:87  */
  assign n9265 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:1050:83  */
  assign n9266 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:1056:87  */
  assign n9267 = is_zero_b & is_inf_a;
  /* TG68K_FPU_ALU.vhd:1056:128  */
  assign n9268 = is_inf_b & is_zero_a;
  /* TG68K_FPU_ALU.vhd:1056:108  */
  assign n9269 = n9267 | n9268;
  /* TG68K_FPU_ALU.vhd:1062:86  */
  assign n9270 = is_inf_a | is_inf_b;
  /* TG68K_FPU_ALU.vhd:1066:87  */
  assign n9271 = is_zero_a | is_zero_b;
  /* TG68K_FPU_ALU.vhd:1072:120  */
  assign n9272 = exp_a + exp_b;
  /* TG68K_FPU_ALU.vhd:1072:138  */
  assign n9274 = n9272 - 15'b011111111111111;
  /* TG68K_FPU_ALU.vhd:1075:82  */
  assign n9275 = mant_a[63:56]; // extract
  /* TG68K_FPU_ALU.vhd:1075:105  */
  assign n9276 = mant_b[63:56]; // extract
  /* TG68K_FPU_ALU.vhd:1075:97  */
  assign n9277 = $unsigned(n9275) > $unsigned(n9276);
  /* TG68K_FPU_ALU.vhd:1075:73  */
  assign n9278 = n9277 ? mant_a : mant_b;
  /* TG68K_FPU_ALU.vhd:1066:65  */
  assign n9280 = n9271 ? 15'b000000000000000 : n9274;
  /* TG68K_FPU_ALU.vhd:1066:65  */
  assign n9282 = n9271 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9278;
  /* TG68K_FPU_ALU.vhd:1066:65  */
  assign n9284 = n9271 ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:1062:65  */
  assign n9286 = n9270 ? 15'b111111111111111 : n9280;
  /* TG68K_FPU_ALU.vhd:1062:65  */
  assign n9288 = n9270 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9282;
  /* TG68K_FPU_ALU.vhd:1062:65  */
  assign n9289 = n9270 ? flags_inexact : n9284;
  /* TG68K_FPU_ALU.vhd:1056:65  */
  assign n9291 = n9269 ? 1'b0 : n9265;
  /* TG68K_FPU_ALU.vhd:1056:65  */
  assign n9293 = n9269 ? 15'b111111111111111 : n9286;
  /* TG68K_FPU_ALU.vhd:1056:65  */
  assign n9295 = n9269 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9288;
  /* TG68K_FPU_ALU.vhd:1056:65  */
  assign n9296 = n9269 ? flags_inexact : n9289;
  /* TG68K_FPU_ALU.vhd:1056:65  */
  assign n9298 = n9269 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:1050:65  */
  assign n9300 = n9266 ? 1'b0 : n9291;
  /* TG68K_FPU_ALU.vhd:1050:65  */
  assign n9302 = n9266 ? 15'b111111111111111 : n9293;
  /* TG68K_FPU_ALU.vhd:1050:65  */
  assign n9304 = n9266 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9295;
  /* TG68K_FPU_ALU.vhd:1050:65  */
  assign n9305 = n9266 ? flags_inexact : n9296;
  /* TG68K_FPU_ALU.vhd:1050:65  */
  assign n9307 = n9266 ? 1'b1 : n9298;
  /* TG68K_FPU_ALU.vhd:1047:57  */
  assign n9309 = operation_code == 7'b0100111;
  /* TG68K_FPU_ALU.vhd:1086:83  */
  assign n9310 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:1086:101  */
  assign n9311 = n9310 | is_inf_a;
  /* TG68K_FPU_ALU.vhd:1086:119  */
  assign n9312 = n9311 | is_zero_b;
  /* TG68K_FPU_ALU.vhd:1100:92  */
  assign n9313 = $unsigned(exp_a) >= $unsigned(exp_b);
  /* TG68K_FPU_ALU.vhd:1105:100  */
  assign n9314 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:1105:118  */
  assign n9316 = $unsigned(n9314) < $unsigned(15'b000000000000111);
  /* TG68K_FPU_ALU.vhd:1108:124  */
  assign n9317 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:1107:129  */
  assign n9319 = n9317[6:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1107:110  */
  assign n9321 = {1'b0, n9319};
  /* TG68K_FPU_ALU.vhd:1111:160  */
  assign n9323 = mant_b + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1111:138  */
  assign n9324 = mant_a % n9323; // umod
  /* TG68K_FPU_ALU.vhd:1112:103  */
  assign n9325 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:1112:121  */
  assign n9327 = $unsigned(n9325) < $unsigned(15'b000000001000000);
  /* TG68K_FPU_ALU.vhd:1116:160  */
  assign n9329 = mant_b + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1116:138  */
  assign n9330 = mant_a % n9329; // umod
  /* TG68K_FPU_ALU.vhd:1112:81  */
  assign n9331 = n9327 ? n9330 : mant_b;
  /* TG68K_FPU_ALU.vhd:1105:81  */
  assign n9332 = n9316 ? n9324 : n9331;
  /* TG68K_FPU_ALU.vhd:1105:81  */
  assign n9334 = n9316 ? n9321 : 8'b01111111;
  /* TG68K_FPU_ALU.vhd:1100:73  */
  assign n9335 = n9313 ? exp_b : exp_a;
  /* TG68K_FPU_ALU.vhd:1100:73  */
  assign n9336 = n9313 ? n9332 : mant_a;
  /* TG68K_FPU_ALU.vhd:1100:73  */
  assign n9338 = n9313 ? n9334 : 8'b00000000;
  /* TG68K_FPU_ALU.vhd:1092:65  */
  assign n9340 = is_zero_a ? 15'b000000000000000 : n9335;
  /* TG68K_FPU_ALU.vhd:1092:65  */
  assign n9342 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9336;
  /* TG68K_FPU_ALU.vhd:1092:65  */
  assign n9343 = is_zero_a ? fmod_quotient : n9338;
  /* TG68K_FPU_ALU.vhd:1092:65  */
  assign n9345 = is_zero_a ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:1086:65  */
  assign n9347 = n9312 ? 1'b0 : sign_a;
  /* TG68K_FPU_ALU.vhd:1086:65  */
  assign n9349 = n9312 ? 15'b111111111111111 : n9340;
  /* TG68K_FPU_ALU.vhd:1086:65  */
  assign n9351 = n9312 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9342;
  /* TG68K_FPU_ALU.vhd:1086:65  */
  assign n9352 = n9312 ? fmod_quotient : n9343;
  /* TG68K_FPU_ALU.vhd:1086:65  */
  assign n9353 = n9312 ? flags_inexact : n9345;
  /* TG68K_FPU_ALU.vhd:1086:65  */
  assign n9355 = n9312 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:1084:57  */
  assign n9357 = operation_code == 7'b0100001;
  /* TG68K_FPU_ALU.vhd:1136:83  */
  assign n9358 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:1136:101  */
  assign n9359 = n9358 | is_inf_a;
  /* TG68K_FPU_ALU.vhd:1136:119  */
  assign n9360 = n9359 | is_zero_b;
  /* TG68K_FPU_ALU.vhd:1150:92  */
  assign n9361 = $unsigned(exp_a) >= $unsigned(exp_b);
  /* TG68K_FPU_ALU.vhd:1153:100  */
  assign n9362 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:1153:118  */
  assign n9364 = $unsigned(n9362) < $unsigned(15'b000000000000111);
  /* TG68K_FPU_ALU.vhd:1156:124  */
  assign n9365 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:1155:129  */
  assign n9367 = n9365[6:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1155:110  */
  assign n9369 = {1'b0, n9367};
  /* TG68K_FPU_ALU.vhd:1159:121  */
  assign n9371 = mant_b >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1161:110  */
  assign n9372 = mant_a[0]; // extract
  /* TG68K_FPU_ALU.vhd:1161:124  */
  assign n9373 = mant_b[0]; // extract
  /* TG68K_FPU_ALU.vhd:1161:114  */
  assign n9374 = n9372 ^ n9373;
  /* TG68K_FPU_ALU.vhd:1162:103  */
  assign n9375 = exp_a - exp_b;
  /* TG68K_FPU_ALU.vhd:1162:121  */
  assign n9377 = $unsigned(n9375) < $unsigned(15'b000000000100000);
  /* TG68K_FPU_ALU.vhd:1166:121  */
  assign n9379 = mant_b >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1167:110  */
  assign n9380 = mant_a[0]; // extract
  /* TG68K_FPU_ALU.vhd:1167:124  */
  assign n9381 = mant_b[0]; // extract
  /* TG68K_FPU_ALU.vhd:1167:114  */
  assign n9382 = n9380 ^ n9381;
  /* TG68K_FPU_ALU.vhd:1171:136  */
  assign n9384 = exp_b - 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:1173:111  */
  assign n9385 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:1162:81  */
  assign n9386 = n9377 ? n9382 : n9385;
  /* TG68K_FPU_ALU.vhd:1162:81  */
  assign n9387 = n9377 ? exp_b : n9384;
  /* TG68K_FPU_ALU.vhd:1162:81  */
  assign n9388 = n9377 ? n9379 : mant_b;
  /* TG68K_FPU_ALU.vhd:1153:81  */
  assign n9389 = n9364 ? n9374 : n9386;
  /* TG68K_FPU_ALU.vhd:1153:81  */
  assign n9390 = n9364 ? exp_b : n9387;
  /* TG68K_FPU_ALU.vhd:1153:81  */
  assign n9391 = n9364 ? n9371 : n9388;
  /* TG68K_FPU_ALU.vhd:1153:81  */
  assign n9393 = n9364 ? n9369 : 8'b01111111;
  /* TG68K_FPU_ALU.vhd:1150:73  */
  assign n9394 = n9361 ? n9389 : sign_a;
  /* TG68K_FPU_ALU.vhd:1150:73  */
  assign n9395 = n9361 ? n9390 : exp_a;
  /* TG68K_FPU_ALU.vhd:1150:73  */
  assign n9396 = n9361 ? n9391 : mant_a;
  /* TG68K_FPU_ALU.vhd:1150:73  */
  assign n9398 = n9361 ? n9393 : 8'b00000000;
  /* TG68K_FPU_ALU.vhd:1142:65  */
  assign n9399 = is_zero_a ? sign_a : n9394;
  /* TG68K_FPU_ALU.vhd:1142:65  */
  assign n9401 = is_zero_a ? 15'b000000000000000 : n9395;
  /* TG68K_FPU_ALU.vhd:1142:65  */
  assign n9403 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9396;
  /* TG68K_FPU_ALU.vhd:1142:65  */
  assign n9404 = is_zero_a ? fmod_quotient : n9398;
  /* TG68K_FPU_ALU.vhd:1142:65  */
  assign n9406 = is_zero_a ? flags_inexact : 1'b1;
  /* TG68K_FPU_ALU.vhd:1136:65  */
  assign n9408 = n9360 ? 1'b0 : n9399;
  /* TG68K_FPU_ALU.vhd:1136:65  */
  assign n9410 = n9360 ? 15'b111111111111111 : n9401;
  /* TG68K_FPU_ALU.vhd:1136:65  */
  assign n9412 = n9360 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9403;
  /* TG68K_FPU_ALU.vhd:1136:65  */
  assign n9413 = n9360 ? fmod_quotient : n9404;
  /* TG68K_FPU_ALU.vhd:1136:65  */
  assign n9414 = n9360 ? flags_inexact : n9406;
  /* TG68K_FPU_ALU.vhd:1136:65  */
  assign n9416 = n9360 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:1134:57  */
  assign n9418 = operation_code == 7'b0100101;
  /* TG68K_FPU_ALU.vhd:1188:83  */
  assign n9419 = is_nan_a | is_nan_b;
  /* TG68K_FPU_ALU.vhd:1206:85  */
  assign n9420 = {16'b0, exp_a};  //  uext
  /* TG68K_FPU_ALU.vhd:1206:73  */
  assign n9421 = {1'b0, n9420};  //  uext
  /* TG68K_FPU_ALU.vhd:1207:82  */
  assign n9423 = $unsigned(exp_b) >= $unsigned(15'b011111111111111);
  /* TG68K_FPU_ALU.vhd:1209:97  */
  assign n9424 = {16'b0, exp_b};  //  uext
  /* TG68K_FPU_ALU.vhd:1209:125  */
  assign n9425 = {1'b0, n9424};  //  uext
  /* TG68K_FPU_ALU.vhd:1209:125  */
  assign n9427 = n9425 - 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:1210:102  */
  assign n9428 = n9421 + n9427;
  /* TG68K_FPU_ALU.vhd:1213:130  */
  assign n9429 = {16'b0, exp_b};  //  uext
  /* TG68K_FPU_ALU.vhd:1213:128  */
  assign n9430 = {1'b0, n9429};  //  uext
  /* TG68K_FPU_ALU.vhd:1213:128  */
  assign n9432 = 32'b00000000000000000011111111111111 - n9430;
  /* TG68K_FPU_ALU.vhd:1214:102  */
  assign n9433 = n9421 - n9432;
  /* TG68K_FPU_ALU.vhd:1207:73  */
  assign n9434 = n9423 ? n9428 : n9433;
  /* TG68K_FPU_ALU.vhd:1218:85  */
  assign n9437 = $signed(n9434) >= $signed(32'b00000000000000000111111111111111);
  /* TG68K_FPU_ALU.vhd:1223:88  */
  assign n9439 = $signed(n9434) <= $signed(32'b00000000000000000000000000000000);
  /* TG68K_FPU_ALU.vhd:1229:124  */
  assign n9440 = n9434[30:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1229:112  */
  assign n9441 = n9440[14:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1223:73  */
  assign n9443 = n9439 ? 15'b000000000000000 : n9441;
  /* TG68K_FPU_ALU.vhd:1223:73  */
  assign n9445 = n9439 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : mant_a;
  /* TG68K_FPU_ALU.vhd:1223:73  */
  assign n9447 = n9439 ? 1'b1 : flags_underflow;
  /* TG68K_FPU_ALU.vhd:1218:73  */
  assign n9449 = n9437 ? 15'b111111111111111 : n9443;
  /* TG68K_FPU_ALU.vhd:1218:73  */
  assign n9451 = n9437 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9445;
  /* TG68K_FPU_ALU.vhd:1218:73  */
  assign n9453 = n9437 ? 1'b1 : flags_overflow;
  /* TG68K_FPU_ALU.vhd:1218:73  */
  assign n9454 = n9437 ? flags_underflow : n9447;
  /* TG68K_FPU_ALU.vhd:1199:65  */
  assign n9456 = is_inf_a ? 15'b111111111111111 : n9449;
  /* TG68K_FPU_ALU.vhd:1199:65  */
  assign n9458 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9451;
  /* TG68K_FPU_ALU.vhd:1199:65  */
  assign n9459 = is_inf_a ? flags_overflow : n9453;
  /* TG68K_FPU_ALU.vhd:1199:65  */
  assign n9460 = is_inf_a ? flags_underflow : n9454;
  /* TG68K_FPU_ALU.vhd:1194:65  */
  assign n9464 = is_zero_a ? 15'b000000000000000 : n9456;
  /* TG68K_FPU_ALU.vhd:1194:65  */
  assign n9466 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9458;
  /* TG68K_FPU_ALU.vhd:1194:65  */
  assign n9467 = is_zero_a ? flags_overflow : n9459;
  /* TG68K_FPU_ALU.vhd:1194:65  */
  assign n9468 = is_zero_a ? flags_underflow : n9460;
  /* TG68K_FPU_ALU.vhd:1188:65  */
  assign n9472 = n9419 ? 1'b0 : sign_a;
  /* TG68K_FPU_ALU.vhd:1188:65  */
  assign n9474 = n9419 ? 15'b111111111111111 : n9464;
  /* TG68K_FPU_ALU.vhd:1188:65  */
  assign n9476 = n9419 ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9466;
  /* TG68K_FPU_ALU.vhd:1188:65  */
  assign n9477 = n9419 ? flags_overflow : n9467;
  /* TG68K_FPU_ALU.vhd:1188:65  */
  assign n9478 = n9419 ? flags_underflow : n9468;
  /* TG68K_FPU_ALU.vhd:1188:65  */
  assign n9480 = n9419 ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:1186:57  */
  assign n9484 = operation_code == 7'b0100110;
  /* TG68K_FPU_ALU.vhd:1254:85  */
  assign n9485 = {16'b0, exp_a};  //  uext
  /* TG68K_FPU_ALU.vhd:1254:113  */
  assign n9486 = {1'b0, n9485};  //  uext
  /* TG68K_FPU_ALU.vhd:1254:113  */
  assign n9488 = n9486 - 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:1256:85  */
  assign n9490 = $signed(n9488) >= $signed(32'b00000000000000000000000000000000);
  /* TG68K_FPU_ALU.vhd:1257:133  */
  assign n9492 = n9488 + 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:1257:124  */
  assign n9493 = n9492[30:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1257:112  */
  assign n9494 = n9493[14:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1260:124  */
  assign n9495 = -n9488;
  /* TG68K_FPU_ALU.vhd:1260:134  */
  assign n9497 = n9495 + 32'b00000000000000000011111111111111;
  /* TG68K_FPU_ALU.vhd:1260:124  */
  assign n9498 = n9497[30:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1260:112  */
  assign n9499 = n9498[14:0];  // trunc
  /* TG68K_FPU_ALU.vhd:1256:73  */
  assign n9502 = n9490 ? 1'b0 : 1'b1;
  /* TG68K_FPU_ALU.vhd:1256:73  */
  assign n9504 = n9490 ? n9494 : n9499;
  /* TG68K_FPU_ALU.vhd:1247:65  */
  assign n9506 = is_zero_a ? 1'b1 : n9502;
  /* TG68K_FPU_ALU.vhd:1247:65  */
  assign n9508 = is_zero_a ? 15'b111111111111111 : n9504;
  /* TG68K_FPU_ALU.vhd:1247:65  */
  assign n9511 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1242:65  */
  assign n9514 = is_inf_a ? 1'b0 : n9506;
  /* TG68K_FPU_ALU.vhd:1242:65  */
  assign n9516 = is_inf_a ? 15'b111111111111111 : n9508;
  /* TG68K_FPU_ALU.vhd:1242:65  */
  assign n9518 = is_inf_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n9511;
  /* TG68K_FPU_ALU.vhd:1237:65  */
  assign n9521 = is_nan_a ? 1'b0 : n9514;
  /* TG68K_FPU_ALU.vhd:1237:65  */
  assign n9523 = is_nan_a ? 15'b111111111111111 : n9516;
  /* TG68K_FPU_ALU.vhd:1237:65  */
  assign n9525 = is_nan_a ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9518;
  /* TG68K_FPU_ALU.vhd:1235:57  */
  assign n9528 = operation_code == 7'b0011110;
  /* TG68K_FPU_ALU.vhd:1279:65  */
  assign n9531 = is_zero_a ? 15'b000000000000000 : 15'b011111111111111;
  /* TG68K_FPU_ALU.vhd:1279:65  */
  assign n9533 = is_zero_a ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : mant_a;
  /* TG68K_FPU_ALU.vhd:1273:65  */
  assign n9535 = is_inf_a ? 1'b0 : sign_a;
  /* TG68K_FPU_ALU.vhd:1273:65  */
  assign n9537 = is_inf_a ? 15'b111111111111111 : n9531;
  /* TG68K_FPU_ALU.vhd:1273:65  */
  assign n9539 = is_inf_a ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9533;
  /* TG68K_FPU_ALU.vhd:1273:65  */
  assign n9541 = is_inf_a ? 1'b1 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:1268:65  */
  assign n9543 = is_nan_a ? 1'b0 : n9535;
  /* TG68K_FPU_ALU.vhd:1268:65  */
  assign n9545 = is_nan_a ? 15'b111111111111111 : n9537;
  /* TG68K_FPU_ALU.vhd:1268:65  */
  assign n9547 = is_nan_a ? 64'b1000000000000000000000000000000000000000000000000000000000000000 : n9539;
  /* TG68K_FPU_ALU.vhd:1268:65  */
  assign n9548 = is_nan_a ? flags_invalid : n9541;
  /* TG68K_FPU_ALU.vhd:1266:57  */
  assign n9550 = operation_code == 7'b0011111;
  assign n9551 = {n9550, n9528, n9484, n9418, n9357, n9309, n9264, n9161, n8675, n8181, n8132, n8018, n7959, n7791, n7601, n7545, n7542, n7540};
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9555 = n9543;
      18'b010000000000000000: n9555 = n9521;
      18'b001000000000000000: n9555 = n9472;
      18'b000100000000000000: n9555 = n9408;
      18'b000010000000000000: n9555 = n9347;
      18'b000001000000000000: n9555 = n9300;
      18'b000000100000000000: n9555 = n9253;
      18'b000000010000000000: n9555 = n9151;
      18'b000000001000000000: n9555 = n8665;
      18'b000000000100000000: n9555 = n8173;
      18'b000000000010000000: n9555 = n8120;
      18'b000000000001000000: n9555 = n8008;
      18'b000000000000100000: n9555 = n7946;
      18'b000000000000010000: n9555 = n7777;
      18'b000000000000001000: n9555 = 1'b0;
      18'b000000000000000100: n9555 = n7543;
      18'b000000000000000010: n9555 = 1'b0;
      18'b000000000000000001: n9555 = sign_b;
      default: n9555 = 1'b0;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9558 = n9545;
      18'b010000000000000000: n9558 = n9523;
      18'b001000000000000000: n9558 = n9474;
      18'b000100000000000000: n9558 = n9410;
      18'b000010000000000000: n9558 = n9349;
      18'b000001000000000000: n9558 = n9302;
      18'b000000100000000000: n9558 = n9255;
      18'b000000010000000000: n9558 = n9153;
      18'b000000001000000000: n9558 = n8667;
      18'b000000000100000000: n9558 = 15'b000000000000000;
      18'b000000000010000000: n9558 = n8122;
      18'b000000000001000000: n9558 = n8010;
      18'b000000000000100000: n9558 = n7948;
      18'b000000000000010000: n9558 = n7779;
      18'b000000000000001000: n9558 = n7593;
      18'b000000000000000100: n9558 = exp_a;
      18'b000000000000000010: n9558 = exp_a;
      18'b000000000000000001: n9558 = exp_b;
      default: n9558 = 15'b000000000000000;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9561 = n9547;
      18'b010000000000000000: n9561 = n9525;
      18'b001000000000000000: n9561 = n9476;
      18'b000100000000000000: n9561 = n9412;
      18'b000010000000000000: n9561 = n9351;
      18'b000001000000000000: n9561 = n9304;
      18'b000000100000000000: n9561 = n9257;
      18'b000000010000000000: n9561 = n9155;
      18'b000000001000000000: n9561 = n8669;
      18'b000000000100000000: n9561 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      18'b000000000010000000: n9561 = n8124;
      18'b000000000001000000: n9561 = n8012;
      18'b000000000000100000: n9561 = n7950;
      18'b000000000000010000: n9561 = n7781;
      18'b000000000000001000: n9561 = n7595;
      18'b000000000000000100: n9561 = mant_a;
      18'b000000000000000010: n9561 = mant_a;
      18'b000000000000000001: n9561 = mant_b;
      default: n9561 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9562 = mant_sum;
      18'b010000000000000000: n9562 = mant_sum;
      18'b001000000000000000: n9562 = mant_sum;
      18'b000100000000000000: n9562 = mant_sum;
      18'b000010000000000000: n9562 = mant_sum;
      18'b000001000000000000: n9562 = mant_sum;
      18'b000000100000000000: n9562 = mant_sum;
      18'b000000010000000000: n9562 = mant_sum;
      18'b000000001000000000: n9562 = mant_sum;
      18'b000000000100000000: n9562 = mant_sum;
      18'b000000000010000000: n9562 = mant_sum;
      18'b000000000001000000: n9562 = mant_sum;
      18'b000000000000100000: n9562 = n7951;
      18'b000000000000010000: n9562 = n7782;
      18'b000000000000001000: n9562 = mant_sum;
      18'b000000000000000100: n9562 = mant_sum;
      18'b000000000000000010: n9562 = mant_sum;
      18'b000000000000000001: n9562 = mant_sum;
      default: n9562 = mant_sum;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9565 = mant_a_aligned;
      18'b010000000000000000: n9565 = mant_a_aligned;
      18'b001000000000000000: n9565 = mant_a_aligned;
      18'b000100000000000000: n9565 = mant_a_aligned;
      18'b000010000000000000: n9565 = mant_a_aligned;
      18'b000001000000000000: n9565 = mant_a_aligned;
      18'b000000100000000000: n9565 = mant_a_aligned;
      18'b000000010000000000: n9565 = mant_a_aligned;
      18'b000000001000000000: n9565 = mant_a_aligned;
      18'b000000000100000000: n9565 = mant_a_aligned;
      18'b000000000010000000: n9565 = mant_a_aligned;
      18'b000000000001000000: n9565 = mant_a_aligned;
      18'b000000000000100000: n9565 = n7953;
      18'b000000000000010000: n9565 = n7785;
      18'b000000000000001000: n9565 = mant_a_aligned;
      18'b000000000000000100: n9565 = mant_a_aligned;
      18'b000000000000000010: n9565 = mant_a_aligned;
      18'b000000000000000001: n9565 = mant_a_aligned;
      default: n9565 = mant_a_aligned;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9566 = mant_b_aligned;
      18'b010000000000000000: n9566 = mant_b_aligned;
      18'b001000000000000000: n9566 = mant_b_aligned;
      18'b000100000000000000: n9566 = mant_b_aligned;
      18'b000010000000000000: n9566 = mant_b_aligned;
      18'b000001000000000000: n9566 = mant_b_aligned;
      18'b000000100000000000: n9566 = mant_b_aligned;
      18'b000000010000000000: n9566 = mant_b_aligned;
      18'b000000001000000000: n9566 = mant_b_aligned;
      18'b000000000100000000: n9566 = mant_b_aligned;
      18'b000000000010000000: n9566 = mant_b_aligned;
      18'b000000000001000000: n9566 = mant_b_aligned;
      18'b000000000000100000: n9566 = n7954;
      18'b000000000000010000: n9566 = n7786;
      18'b000000000000001000: n9566 = mant_b_aligned;
      18'b000000000000000100: n9566 = mant_b_aligned;
      18'b000000000000000010: n9566 = mant_b_aligned;
      18'b000000000000000001: n9566 = mant_b_aligned;
      default: n9566 = mant_b_aligned;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9567 = exp_larger;
      18'b010000000000000000: n9567 = exp_larger;
      18'b001000000000000000: n9567 = exp_larger;
      18'b000100000000000000: n9567 = exp_larger;
      18'b000010000000000000: n9567 = exp_larger;
      18'b000001000000000000: n9567 = exp_larger;
      18'b000000100000000000: n9567 = exp_larger;
      18'b000000010000000000: n9567 = exp_larger;
      18'b000000001000000000: n9567 = exp_larger;
      18'b000000000100000000: n9567 = exp_larger;
      18'b000000000010000000: n9567 = exp_larger;
      18'b000000000001000000: n9567 = exp_larger;
      18'b000000000000100000: n9567 = n7955;
      18'b000000000000010000: n9567 = n7787;
      18'b000000000000001000: n9567 = exp_larger;
      18'b000000000000000100: n9567 = exp_larger;
      18'b000000000000000010: n9567 = exp_larger;
      18'b000000000000000001: n9567 = exp_larger;
      default: n9567 = exp_larger;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9569 = mult_result;
      18'b010000000000000000: n9569 = mult_result;
      18'b001000000000000000: n9569 = mult_result;
      18'b000100000000000000: n9569 = mult_result;
      18'b000010000000000000: n9569 = mult_result;
      18'b000001000000000000: n9569 = mult_result;
      18'b000000100000000000: n9569 = mult_result;
      18'b000000010000000000: n9569 = mult_result;
      18'b000000001000000000: n9569 = mult_result;
      18'b000000000100000000: n9569 = mult_result;
      18'b000000000010000000: n9569 = mult_result;
      18'b000000000001000000: n9569 = n8013;
      18'b000000000000100000: n9569 = mult_result;
      18'b000000000000010000: n9569 = mult_result;
      18'b000000000000001000: n9569 = mult_result;
      18'b000000000000000100: n9569 = mult_result;
      18'b000000000000000010: n9569 = mult_result;
      18'b000000000000000001: n9569 = mult_result;
      default: n9569 = mult_result;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9570 = fmod_quotient;
      18'b010000000000000000: n9570 = fmod_quotient;
      18'b001000000000000000: n9570 = fmod_quotient;
      18'b000100000000000000: n9570 = n9413;
      18'b000010000000000000: n9570 = n9352;
      18'b000001000000000000: n9570 = fmod_quotient;
      18'b000000100000000000: n9570 = fmod_quotient;
      18'b000000010000000000: n9570 = fmod_quotient;
      18'b000000001000000000: n9570 = fmod_quotient;
      18'b000000000100000000: n9570 = fmod_quotient;
      18'b000000000010000000: n9570 = fmod_quotient;
      18'b000000000001000000: n9570 = fmod_quotient;
      18'b000000000000100000: n9570 = fmod_quotient;
      18'b000000000000010000: n9570 = fmod_quotient;
      18'b000000000000001000: n9570 = fmod_quotient;
      18'b000000000000000100: n9570 = fmod_quotient;
      18'b000000000000000010: n9570 = fmod_quotient;
      18'b000000000000000001: n9570 = fmod_quotient;
      default: n9570 = fmod_quotient;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9571 = flags_overflow;
      18'b010000000000000000: n9571 = flags_overflow;
      18'b001000000000000000: n9571 = n9477;
      18'b000100000000000000: n9571 = flags_overflow;
      18'b000010000000000000: n9571 = flags_overflow;
      18'b000001000000000000: n9571 = flags_overflow;
      18'b000000100000000000: n9571 = n9258;
      18'b000000010000000000: n9571 = flags_overflow;
      18'b000000001000000000: n9571 = flags_overflow;
      18'b000000000100000000: n9571 = flags_overflow;
      18'b000000000010000000: n9571 = n8126;
      18'b000000000001000000: n9571 = flags_overflow;
      18'b000000000000100000: n9571 = flags_overflow;
      18'b000000000000010000: n9571 = flags_overflow;
      18'b000000000000001000: n9571 = flags_overflow;
      18'b000000000000000100: n9571 = flags_overflow;
      18'b000000000000000010: n9571 = flags_overflow;
      18'b000000000000000001: n9571 = flags_overflow;
      default: n9571 = flags_overflow;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9572 = flags_underflow;
      18'b010000000000000000: n9572 = flags_underflow;
      18'b001000000000000000: n9572 = n9478;
      18'b000100000000000000: n9572 = flags_underflow;
      18'b000010000000000000: n9572 = flags_underflow;
      18'b000001000000000000: n9572 = flags_underflow;
      18'b000000100000000000: n9572 = flags_underflow;
      18'b000000010000000000: n9572 = flags_underflow;
      18'b000000001000000000: n9572 = flags_underflow;
      18'b000000000100000000: n9572 = flags_underflow;
      18'b000000000010000000: n9572 = flags_underflow;
      18'b000000000001000000: n9572 = flags_underflow;
      18'b000000000000100000: n9572 = flags_underflow;
      18'b000000000000010000: n9572 = flags_underflow;
      18'b000000000000001000: n9572 = flags_underflow;
      18'b000000000000000100: n9572 = flags_underflow;
      18'b000000000000000010: n9572 = flags_underflow;
      18'b000000000000000001: n9572 = flags_underflow;
      default: n9572 = flags_underflow;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9573 = flags_inexact;
      18'b010000000000000000: n9573 = flags_inexact;
      18'b001000000000000000: n9573 = flags_inexact;
      18'b000100000000000000: n9573 = n9414;
      18'b000010000000000000: n9573 = n9353;
      18'b000001000000000000: n9573 = n9305;
      18'b000000100000000000: n9573 = n9259;
      18'b000000010000000000: n9573 = n9156;
      18'b000000001000000000: n9573 = n8670;
      18'b000000000100000000: n9573 = flags_inexact;
      18'b000000000010000000: n9573 = n8127;
      18'b000000000001000000: n9573 = n8014;
      18'b000000000000100000: n9573 = flags_inexact;
      18'b000000000000010000: n9573 = flags_inexact;
      18'b000000000000001000: n9573 = n7596;
      18'b000000000000000100: n9573 = flags_inexact;
      18'b000000000000000010: n9573 = flags_inexact;
      18'b000000000000000001: n9573 = flags_inexact;
      default: n9573 = flags_inexact;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9575 = n9548;
      18'b010000000000000000: n9575 = flags_invalid;
      18'b001000000000000000: n9575 = n9480;
      18'b000100000000000000: n9575 = n9416;
      18'b000010000000000000: n9575 = n9355;
      18'b000001000000000000: n9575 = n9307;
      18'b000000100000000000: n9575 = n9261;
      18'b000000010000000000: n9575 = n9158;
      18'b000000001000000000: n9575 = n8672;
      18'b000000000100000000: n9575 = n8176;
      18'b000000000010000000: n9575 = n8129;
      18'b000000000001000000: n9575 = n8016;
      18'b000000000000100000: n9575 = n7957;
      18'b000000000000010000: n9575 = n7789;
      18'b000000000000001000: n9575 = n7598;
      18'b000000000000000100: n9575 = flags_invalid;
      18'b000000000000000010: n9575 = flags_invalid;
      18'b000000000000000001: n9575 = flags_invalid;
      default: n9575 = 1'b1;
    endcase
  /* TG68K_FPU_ALU.vhd:339:49  */
  always @*
    case (n9551)
      18'b100000000000000000: n9576 = flags_div_by_zero;
      18'b010000000000000000: n9576 = flags_div_by_zero;
      18'b001000000000000000: n9576 = flags_div_by_zero;
      18'b000100000000000000: n9576 = flags_div_by_zero;
      18'b000010000000000000: n9576 = flags_div_by_zero;
      18'b000001000000000000: n9576 = flags_div_by_zero;
      18'b000000100000000000: n9576 = n9262;
      18'b000000010000000000: n9576 = flags_div_by_zero;
      18'b000000001000000000: n9576 = flags_div_by_zero;
      18'b000000000100000000: n9576 = flags_div_by_zero;
      18'b000000000010000000: n9576 = n8130;
      18'b000000000001000000: n9576 = flags_div_by_zero;
      18'b000000000000100000: n9576 = flags_div_by_zero;
      18'b000000000000010000: n9576 = flags_div_by_zero;
      18'b000000000000001000: n9576 = flags_div_by_zero;
      18'b000000000000000100: n9576 = flags_div_by_zero;
      18'b000000000000000010: n9576 = flags_div_by_zero;
      18'b000000000000000001: n9576 = flags_div_by_zero;
      default: n9576 = flags_div_by_zero;
    endcase
  /* TG68K_FPU_ALU.vhd:338:41  */
  assign n9580 = alu_state == 3'b011;
  /* TG68K_FPU_ALU.vhd:1304:63  */
  assign n9582 = exp_result == 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:1304:89  */
  assign n9584 = mant_result == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1304:74  */
  assign n9585 = n9582 | n9584;
  /* TG68K_FPU_ALU.vhd:1308:66  */
  assign n9587 = $unsigned(exp_result) >= $unsigned(15'b111111111111111);
  /* TG68K_FPU_ALU.vhd:1313:65  */
  assign n9588 = exp_result[14]; // extract
  /* TG68K_FPU_ALU.vhd:1321:71  */
  assign n9589 = mant_result[63]; // extract
  /* TG68K_FPU_ALU.vhd:1321:76  */
  assign n9590 = ~n9589;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9592 = mant_result[63]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9598 = n9592 ? 1'b0 : 1'b1;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9600 = mant_result[62]; // extract
  /* TG68K_FPU_ALU.vhd:1327:81  */
  assign n9603 = n9598 ? 6'b000001 : 6'b000000;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9607 = n9616 ? 1'b0 : n9598;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9610 = n9600 ? n9603 : 6'b000000;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9611 = n9598 & n9600;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9614 = n9598 ? n9610 : 6'b000000;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9616 = n9611 & n9598;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9617 = mant_result[61]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9619 = n9628 ? 6'b000010 : n9614;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9623 = n9629 ? 1'b0 : n9607;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9625 = n9607 & n9617;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9626 = n9607 & n9617;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9628 = n9625 & n9607;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9629 = n9626 & n9607;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9630 = mant_result[60]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9632 = n9641 ? 6'b000011 : n9619;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9636 = n9642 ? 1'b0 : n9623;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9638 = n9623 & n9630;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9639 = n9623 & n9630;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9641 = n9638 & n9623;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9642 = n9639 & n9623;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9643 = mant_result[59]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9645 = n9654 ? 6'b000100 : n9632;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9649 = n9655 ? 1'b0 : n9636;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9651 = n9636 & n9643;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9652 = n9636 & n9643;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9654 = n9651 & n9636;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9655 = n9652 & n9636;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9656 = mant_result[58]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9658 = n9667 ? 6'b000101 : n9645;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9662 = n9668 ? 1'b0 : n9649;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9664 = n9649 & n9656;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9665 = n9649 & n9656;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9667 = n9664 & n9649;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9668 = n9665 & n9649;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9669 = mant_result[57]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9671 = n9680 ? 6'b000110 : n9658;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9675 = n9681 ? 1'b0 : n9662;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9677 = n9662 & n9669;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9678 = n9662 & n9669;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9680 = n9677 & n9662;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9681 = n9678 & n9662;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9682 = mant_result[56]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9684 = n9693 ? 6'b000111 : n9671;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9688 = n9694 ? 1'b0 : n9675;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9690 = n9675 & n9682;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9691 = n9675 & n9682;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9693 = n9690 & n9675;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9694 = n9691 & n9675;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9695 = mant_result[55]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9697 = n9706 ? 6'b001000 : n9684;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9701 = n9707 ? 1'b0 : n9688;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9703 = n9688 & n9695;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9704 = n9688 & n9695;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9706 = n9703 & n9688;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9707 = n9704 & n9688;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9708 = mant_result[54]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9710 = n9719 ? 6'b001001 : n9697;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9714 = n9720 ? 1'b0 : n9701;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9716 = n9701 & n9708;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9717 = n9701 & n9708;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9719 = n9716 & n9701;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9720 = n9717 & n9701;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9721 = mant_result[53]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9723 = n9732 ? 6'b001010 : n9710;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9727 = n9733 ? 1'b0 : n9714;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9729 = n9714 & n9721;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9730 = n9714 & n9721;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9732 = n9729 & n9714;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9733 = n9730 & n9714;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9734 = mant_result[52]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9736 = n9745 ? 6'b001011 : n9723;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9740 = n9746 ? 1'b0 : n9727;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9742 = n9727 & n9734;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9743 = n9727 & n9734;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9745 = n9742 & n9727;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9746 = n9743 & n9727;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9747 = mant_result[51]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9749 = n9758 ? 6'b001100 : n9736;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9753 = n9759 ? 1'b0 : n9740;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9755 = n9740 & n9747;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9756 = n9740 & n9747;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9758 = n9755 & n9740;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9759 = n9756 & n9740;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9760 = mant_result[50]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9762 = n9771 ? 6'b001101 : n9749;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9766 = n9772 ? 1'b0 : n9753;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9768 = n9753 & n9760;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9769 = n9753 & n9760;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9771 = n9768 & n9753;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9772 = n9769 & n9753;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9773 = mant_result[49]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9775 = n9784 ? 6'b001110 : n9762;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9779 = n9785 ? 1'b0 : n9766;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9781 = n9766 & n9773;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9782 = n9766 & n9773;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9784 = n9781 & n9766;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9785 = n9782 & n9766;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9786 = mant_result[48]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9788 = n9797 ? 6'b001111 : n9775;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9792 = n9798 ? 1'b0 : n9779;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9794 = n9779 & n9786;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9795 = n9779 & n9786;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9797 = n9794 & n9779;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9798 = n9795 & n9779;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9799 = mant_result[47]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9801 = n9810 ? 6'b010000 : n9788;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9805 = n9811 ? 1'b0 : n9792;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9807 = n9792 & n9799;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9808 = n9792 & n9799;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9810 = n9807 & n9792;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9811 = n9808 & n9792;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9812 = mant_result[46]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9814 = n9823 ? 6'b010001 : n9801;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9818 = n9824 ? 1'b0 : n9805;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9820 = n9805 & n9812;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9821 = n9805 & n9812;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9823 = n9820 & n9805;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9824 = n9821 & n9805;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9825 = mant_result[45]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9827 = n9836 ? 6'b010010 : n9814;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9831 = n9837 ? 1'b0 : n9818;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9833 = n9818 & n9825;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9834 = n9818 & n9825;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9836 = n9833 & n9818;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9837 = n9834 & n9818;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9838 = mant_result[44]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9840 = n9849 ? 6'b010011 : n9827;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9844 = n9850 ? 1'b0 : n9831;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9846 = n9831 & n9838;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9847 = n9831 & n9838;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9849 = n9846 & n9831;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9850 = n9847 & n9831;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9851 = mant_result[43]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9853 = n9862 ? 6'b010100 : n9840;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9857 = n9863 ? 1'b0 : n9844;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9859 = n9844 & n9851;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9860 = n9844 & n9851;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9862 = n9859 & n9844;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9863 = n9860 & n9844;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9864 = mant_result[42]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9866 = n9875 ? 6'b010101 : n9853;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9870 = n9876 ? 1'b0 : n9857;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9872 = n9857 & n9864;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9873 = n9857 & n9864;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9875 = n9872 & n9857;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9876 = n9873 & n9857;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9877 = mant_result[41]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9879 = n9888 ? 6'b010110 : n9866;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9883 = n9889 ? 1'b0 : n9870;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9885 = n9870 & n9877;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9886 = n9870 & n9877;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9888 = n9885 & n9870;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9889 = n9886 & n9870;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9890 = mant_result[40]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9892 = n9901 ? 6'b010111 : n9879;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9896 = n9902 ? 1'b0 : n9883;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9898 = n9883 & n9890;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9899 = n9883 & n9890;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9901 = n9898 & n9883;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9902 = n9899 & n9883;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9903 = mant_result[39]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9905 = n9914 ? 6'b011000 : n9892;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9909 = n9915 ? 1'b0 : n9896;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9911 = n9896 & n9903;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9912 = n9896 & n9903;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9914 = n9911 & n9896;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9915 = n9912 & n9896;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9916 = mant_result[38]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9918 = n9927 ? 6'b011001 : n9905;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9922 = n9928 ? 1'b0 : n9909;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9924 = n9909 & n9916;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9925 = n9909 & n9916;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9927 = n9924 & n9909;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9928 = n9925 & n9909;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9929 = mant_result[37]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9931 = n9940 ? 6'b011010 : n9918;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9935 = n9941 ? 1'b0 : n9922;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9937 = n9922 & n9929;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9938 = n9922 & n9929;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9940 = n9937 & n9922;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9941 = n9938 & n9922;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9942 = mant_result[36]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9944 = n9953 ? 6'b011011 : n9931;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9948 = n9954 ? 1'b0 : n9935;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9950 = n9935 & n9942;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9951 = n9935 & n9942;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9953 = n9950 & n9935;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9954 = n9951 & n9935;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9955 = mant_result[35]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9957 = n9966 ? 6'b011100 : n9944;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9961 = n9967 ? 1'b0 : n9948;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9963 = n9948 & n9955;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9964 = n9948 & n9955;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9966 = n9963 & n9948;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9967 = n9964 & n9948;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9968 = mant_result[34]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9970 = n9979 ? 6'b011101 : n9957;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9974 = n9980 ? 1'b0 : n9961;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9976 = n9961 & n9968;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9977 = n9961 & n9968;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9979 = n9976 & n9961;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9980 = n9977 & n9961;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9981 = mant_result[33]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9983 = n9992 ? 6'b011110 : n9970;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9987 = n9993 ? 1'b0 : n9974;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9989 = n9974 & n9981;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9990 = n9974 & n9981;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9992 = n9989 & n9974;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9993 = n9990 & n9974;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n9994 = mant_result[32]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n9996 = n10005 ? 6'b011111 : n9983;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10000 = n10006 ? 1'b0 : n9987;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10002 = n9987 & n9994;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10003 = n9987 & n9994;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10005 = n10002 & n9987;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10006 = n10003 & n9987;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10007 = mant_result[31]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10009 = n10018 ? 6'b100000 : n9996;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10013 = n10019 ? 1'b0 : n10000;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10015 = n10000 & n10007;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10016 = n10000 & n10007;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10018 = n10015 & n10000;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10019 = n10016 & n10000;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10020 = mant_result[30]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10022 = n10031 ? 6'b100001 : n10009;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10026 = n10032 ? 1'b0 : n10013;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10028 = n10013 & n10020;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10029 = n10013 & n10020;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10031 = n10028 & n10013;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10032 = n10029 & n10013;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10033 = mant_result[29]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10035 = n10044 ? 6'b100010 : n10022;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10039 = n10045 ? 1'b0 : n10026;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10041 = n10026 & n10033;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10042 = n10026 & n10033;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10044 = n10041 & n10026;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10045 = n10042 & n10026;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10046 = mant_result[28]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10048 = n10057 ? 6'b100011 : n10035;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10052 = n10058 ? 1'b0 : n10039;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10054 = n10039 & n10046;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10055 = n10039 & n10046;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10057 = n10054 & n10039;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10058 = n10055 & n10039;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10059 = mant_result[27]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10061 = n10070 ? 6'b100100 : n10048;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10065 = n10071 ? 1'b0 : n10052;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10067 = n10052 & n10059;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10068 = n10052 & n10059;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10070 = n10067 & n10052;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10071 = n10068 & n10052;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10072 = mant_result[26]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10074 = n10083 ? 6'b100101 : n10061;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10078 = n10084 ? 1'b0 : n10065;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10080 = n10065 & n10072;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10081 = n10065 & n10072;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10083 = n10080 & n10065;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10084 = n10081 & n10065;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10085 = mant_result[25]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10087 = n10096 ? 6'b100110 : n10074;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10091 = n10097 ? 1'b0 : n10078;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10093 = n10078 & n10085;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10094 = n10078 & n10085;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10096 = n10093 & n10078;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10097 = n10094 & n10078;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10098 = mant_result[24]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10100 = n10109 ? 6'b100111 : n10087;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10104 = n10110 ? 1'b0 : n10091;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10106 = n10091 & n10098;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10107 = n10091 & n10098;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10109 = n10106 & n10091;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10110 = n10107 & n10091;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10111 = mant_result[23]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10113 = n10122 ? 6'b101000 : n10100;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10117 = n10123 ? 1'b0 : n10104;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10119 = n10104 & n10111;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10120 = n10104 & n10111;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10122 = n10119 & n10104;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10123 = n10120 & n10104;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10124 = mant_result[22]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10126 = n10135 ? 6'b101001 : n10113;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10130 = n10136 ? 1'b0 : n10117;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10132 = n10117 & n10124;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10133 = n10117 & n10124;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10135 = n10132 & n10117;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10136 = n10133 & n10117;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10137 = mant_result[21]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10139 = n10148 ? 6'b101010 : n10126;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10143 = n10149 ? 1'b0 : n10130;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10145 = n10130 & n10137;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10146 = n10130 & n10137;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10148 = n10145 & n10130;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10149 = n10146 & n10130;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10150 = mant_result[20]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10152 = n10161 ? 6'b101011 : n10139;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10156 = n10162 ? 1'b0 : n10143;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10158 = n10143 & n10150;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10159 = n10143 & n10150;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10161 = n10158 & n10143;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10162 = n10159 & n10143;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10163 = mant_result[19]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10165 = n10174 ? 6'b101100 : n10152;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10169 = n10175 ? 1'b0 : n10156;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10171 = n10156 & n10163;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10172 = n10156 & n10163;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10174 = n10171 & n10156;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10175 = n10172 & n10156;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10176 = mant_result[18]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10178 = n10187 ? 6'b101101 : n10165;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10182 = n10188 ? 1'b0 : n10169;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10184 = n10169 & n10176;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10185 = n10169 & n10176;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10187 = n10184 & n10169;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10188 = n10185 & n10169;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10189 = mant_result[17]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10191 = n10200 ? 6'b101110 : n10178;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10195 = n10201 ? 1'b0 : n10182;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10197 = n10182 & n10189;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10198 = n10182 & n10189;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10200 = n10197 & n10182;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10201 = n10198 & n10182;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10202 = mant_result[16]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10204 = n10213 ? 6'b101111 : n10191;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10208 = n10214 ? 1'b0 : n10195;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10210 = n10195 & n10202;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10211 = n10195 & n10202;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10213 = n10210 & n10195;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10214 = n10211 & n10195;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10215 = mant_result[15]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10217 = n10226 ? 6'b110000 : n10204;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10221 = n10227 ? 1'b0 : n10208;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10223 = n10208 & n10215;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10224 = n10208 & n10215;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10226 = n10223 & n10208;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10227 = n10224 & n10208;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10228 = mant_result[14]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10230 = n10239 ? 6'b110001 : n10217;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10234 = n10240 ? 1'b0 : n10221;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10236 = n10221 & n10228;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10237 = n10221 & n10228;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10239 = n10236 & n10221;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10240 = n10237 & n10221;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10241 = mant_result[13]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10243 = n10252 ? 6'b110010 : n10230;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10247 = n10253 ? 1'b0 : n10234;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10249 = n10234 & n10241;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10250 = n10234 & n10241;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10252 = n10249 & n10234;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10253 = n10250 & n10234;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10254 = mant_result[12]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10256 = n10265 ? 6'b110011 : n10243;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10260 = n10266 ? 1'b0 : n10247;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10262 = n10247 & n10254;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10263 = n10247 & n10254;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10265 = n10262 & n10247;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10266 = n10263 & n10247;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10267 = mant_result[11]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10269 = n10278 ? 6'b110100 : n10256;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10273 = n10279 ? 1'b0 : n10260;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10275 = n10260 & n10267;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10276 = n10260 & n10267;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10278 = n10275 & n10260;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10279 = n10276 & n10260;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10280 = mant_result[10]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10282 = n10291 ? 6'b110101 : n10269;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10286 = n10292 ? 1'b0 : n10273;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10288 = n10273 & n10280;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10289 = n10273 & n10280;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10291 = n10288 & n10273;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10292 = n10289 & n10273;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10293 = mant_result[9]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10295 = n10304 ? 6'b110110 : n10282;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10299 = n10305 ? 1'b0 : n10286;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10301 = n10286 & n10293;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10302 = n10286 & n10293;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10304 = n10301 & n10286;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10305 = n10302 & n10286;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10306 = mant_result[8]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10308 = n10317 ? 6'b110111 : n10295;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10312 = n10318 ? 1'b0 : n10299;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10314 = n10299 & n10306;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10315 = n10299 & n10306;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10317 = n10314 & n10299;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10318 = n10315 & n10299;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10319 = mant_result[7]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10321 = n10330 ? 6'b111000 : n10308;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10325 = n10331 ? 1'b0 : n10312;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10327 = n10312 & n10319;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10328 = n10312 & n10319;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10330 = n10327 & n10312;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10331 = n10328 & n10312;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10332 = mant_result[6]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10334 = n10343 ? 6'b111001 : n10321;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10338 = n10344 ? 1'b0 : n10325;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10340 = n10325 & n10332;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10341 = n10325 & n10332;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10343 = n10340 & n10325;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10344 = n10341 & n10325;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10345 = mant_result[5]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10347 = n10356 ? 6'b111010 : n10334;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10351 = n10357 ? 1'b0 : n10338;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10353 = n10338 & n10345;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10354 = n10338 & n10345;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10356 = n10353 & n10338;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10357 = n10354 & n10338;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10358 = mant_result[4]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10360 = n10369 ? 6'b111011 : n10347;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10364 = n10370 ? 1'b0 : n10351;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10366 = n10351 & n10358;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10367 = n10351 & n10358;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10369 = n10366 & n10351;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10370 = n10367 & n10351;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10371 = mant_result[3]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10373 = n10382 ? 6'b111100 : n10360;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10377 = n10383 ? 1'b0 : n10364;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10379 = n10364 & n10371;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10380 = n10364 & n10371;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10382 = n10379 & n10364;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10383 = n10380 & n10364;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10384 = mant_result[2]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10386 = n10395 ? 6'b111101 : n10373;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10390 = n10396 ? 1'b0 : n10377;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10392 = n10377 & n10384;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10393 = n10377 & n10384;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10395 = n10392 & n10377;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10396 = n10393 & n10377;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10397 = mant_result[1]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10399 = n10408 ? 6'b111110 : n10386;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10403 = n10409 ? 1'b0 : n10390;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10405 = n10390 & n10397;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10406 = n10390 & n10397;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10408 = n10405 & n10390;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10409 = n10406 & n10390;
  /* TG68K_FPU_ALU.vhd:1326:87  */
  assign n10410 = mant_result[0]; // extract
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10412 = n10421 ? 6'b111111 : n10399;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10418 = n10403 & n10410;
  /* TG68K_FPU_ALU.vhd:1326:73  */
  assign n10421 = n10418 & n10403;
  /* TG68K_FPU_ALU.vhd:1333:79  */
  assign n10423 = {26'b0, n10412};  //  uext
  /* TG68K_FPU_ALU.vhd:1333:79  */
  assign n10425 = n10423 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1333:99  */
  assign n10427 = mant_result == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1333:83  */
  assign n10428 = n10427 & n10425;
  /* TG68K_FPU_ALU.vhd:1342:99  */
  assign n10429 = sign_a == sign_b;
  /* TG68K_FPU_ALU.vhd:1344:109  */
  assign n10431 = rounding_mode == 2'b11;
  /* TG68K_FPU_ALU.vhd:1344:89  */
  assign n10434 = n10431 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1342:89  */
  assign n10435 = n10429 ? sign_a : n10434;
  /* TG68K_FPU_ALU.vhd:1340:81  */
  assign n10437 = operation_code == 7'b0100010;
  /* TG68K_FPU_ALU.vhd:1351:99  */
  assign n10438 = ~sign_a;
  /* TG68K_FPU_ALU.vhd:1351:116  */
  assign n10439 = ~sign_b;
  /* TG68K_FPU_ALU.vhd:1351:105  */
  assign n10440 = n10439 & n10438;
  /* TG68K_FPU_ALU.vhd:1353:108  */
  assign n10441 = sign_b & sign_a;
  /* TG68K_FPU_ALU.vhd:1355:102  */
  assign n10442 = ~sign_a;
  /* TG68K_FPU_ALU.vhd:1355:108  */
  assign n10443 = sign_b & n10442;
  /* TG68K_FPU_ALU.vhd:1355:89  */
  assign n10446 = n10443 ? 1'b0 : 1'b1;
  /* TG68K_FPU_ALU.vhd:1353:89  */
  assign n10448 = n10441 ? 1'b0 : n10446;
  /* TG68K_FPU_ALU.vhd:1351:89  */
  assign n10450 = n10440 ? 1'b0 : n10448;
  /* TG68K_FPU_ALU.vhd:1349:81  */
  assign n10452 = operation_code == 7'b0101000;
  /* TG68K_FPU_ALU.vhd:1362:111  */
  assign n10453 = sign_a ^ sign_b;
  /* TG68K_FPU_ALU.vhd:1360:81  */
  assign n10455 = operation_code == 7'b0100011;
  /* TG68K_FPU_ALU.vhd:1360:94  */
  assign n10457 = operation_code == 7'b0100000;
  /* TG68K_FPU_ALU.vhd:1360:94  */
  assign n10458 = n10455 | n10457;
  /* TG68K_FPU_ALU.vhd:1360:104  */
  assign n10460 = operation_code == 7'b0100100;
  /* TG68K_FPU_ALU.vhd:1360:104  */
  assign n10461 = n10458 | n10460;
  assign n10462 = {n10461, n10452, n10437};
  /* TG68K_FPU_ALU.vhd:1339:73  */
  always @*
    case (n10462)
      3'b100: n10463 = n10453;
      3'b010: n10463 = n10450;
      3'b001: n10463 = n10435;
      default: n10463 = sign_result;
    endcase
  /* TG68K_FPU_ALU.vhd:1368:82  */
  assign n10464 = {26'b0, n10412};  //  uext
  /* TG68K_FPU_ALU.vhd:1368:82  */
  assign n10466 = $signed(n10464) > $signed(32'b00000000000000000000000000000000);
  /* TG68K_FPU_ALU.vhd:1368:101  */
  assign n10467 = {26'b0, n10412};  //  uext
  /* TG68K_FPU_ALU.vhd:1368:101  */
  assign n10469 = $signed(n10467) <= $signed(32'b00000000000000000000000000111111);
  /* TG68K_FPU_ALU.vhd:1368:86  */
  assign n10470 = n10469 & n10466;
  /* TG68K_FPU_ALU.vhd:1369:76  */
  assign n10471 = {16'b0, exp_result};  //  uext
  /* TG68K_FPU_ALU.vhd:1369:109  */
  assign n10472 = {1'b0, n10471};  //  uext
  /* TG68K_FPU_ALU.vhd:1369:109  */
  assign n10473 = {26'b0, n10412};  //  uext
  /* TG68K_FPU_ALU.vhd:1369:109  */
  assign n10474 = $signed(n10472) > $signed(n10473);
  /* TG68K_FPU_ALU.vhd:1371:135  */
  assign n10476 = {9'b0, n10412};  //  uext
  /* TG68K_FPU_ALU.vhd:1371:133  */
  assign n10477 = exp_result - n10476;
  /* TG68K_FPU_ALU.vhd:1372:147  */
  assign n10478 = {25'b0, n10412};  //  uext
  /* TG68K_FPU_ALU.vhd:1372:113  */
  assign n10479 = mant_result << n10478;
  /* TG68K_FPU_ALU.vhd:1379:95  */
  assign n10480 = mant_result[63]; // extract
  /* TG68K_FPU_ALU.vhd:1381:121  */
  assign n10482 = mant_result >> 31'b0000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1379:81  */
  assign n10484 = n10480 ? n10482 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1369:73  */
  assign n10486 = n10474 ? n10477 : 15'b000000000000000;
  /* TG68K_FPU_ALU.vhd:1369:73  */
  assign n10487 = n10474 ? n10479 : n10484;
  /* TG68K_FPU_ALU.vhd:1369:73  */
  assign n10489 = n10474 ? flags_underflow : 1'b1;
  /* TG68K_FPU_ALU.vhd:1368:65  */
  assign n10490 = n10470 ? n10486 : exp_result;
  /* TG68K_FPU_ALU.vhd:1368:65  */
  assign n10491 = n10470 ? n10487 : mant_result;
  /* TG68K_FPU_ALU.vhd:1368:65  */
  assign n10492 = n10470 ? n10489 : flags_underflow;
  /* TG68K_FPU_ALU.vhd:1321:57  */
  assign n10493 = n10500 ? n10463 : sign_result;
  /* TG68K_FPU_ALU.vhd:1333:65  */
  assign n10495 = n10428 ? 15'b000000000000000 : n10490;
  /* TG68K_FPU_ALU.vhd:1333:65  */
  assign n10497 = n10428 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n10491;
  /* TG68K_FPU_ALU.vhd:1333:65  */
  assign n10499 = n10428 ? 1'b1 : n10492;
  /* TG68K_FPU_ALU.vhd:1321:57  */
  assign n10500 = n10428 & n9590;
  /* TG68K_FPU_ALU.vhd:1321:57  */
  assign n10501 = n9590 ? n10495 : exp_result;
  /* TG68K_FPU_ALU.vhd:1321:57  */
  assign n10502 = n9590 ? n10497 : mant_result;
  /* TG68K_FPU_ALU.vhd:1321:57  */
  assign n10503 = n9590 ? n10499 : flags_underflow;
  /* TG68K_FPU_ALU.vhd:1399:84  */
  assign n10505 = mant_sum[64]; // extract
  /* TG68K_FPU_ALU.vhd:1401:102  */
  assign n10506 = mant_sum[1]; // extract
  /* TG68K_FPU_ALU.vhd:1402:102  */
  assign n10507 = mant_sum[0]; // extract
  /* TG68K_FPU_ALU.vhd:1406:102  */
  assign n10508 = mant_sum[0]; // extract
  /* TG68K_FPU_ALU.vhd:1399:73  */
  assign n10509 = n10505 ? n10506 : n10508;
  /* TG68K_FPU_ALU.vhd:1399:73  */
  assign n10511 = n10505 ? n10507 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1397:65  */
  assign n10513 = operation_code == 7'b0100010;
  /* TG68K_FPU_ALU.vhd:1397:78  */
  assign n10515 = operation_code == 7'b0101000;
  /* TG68K_FPU_ALU.vhd:1397:78  */
  assign n10516 = n10513 | n10515;
  /* TG68K_FPU_ALU.vhd:1412:97  */
  assign n10517 = mult_result[63]; // extract
  /* TG68K_FPU_ALU.vhd:1413:97  */
  assign n10518 = mult_result[62]; // extract
  /* TG68K_FPU_ALU.vhd:1415:87  */
  assign n10519 = mult_result[61:0]; // extract
  /* TG68K_FPU_ALU.vhd:1415:101  */
  assign n10521 = n10519 != 62'b00000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1415:73  */
  assign n10524 = n10521 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1410:65  */
  assign n10526 = operation_code == 7'b0100011;
  /* TG68K_FPU_ALU.vhd:1425:97  */
  assign n10527 = mant_result[0]; // extract
  /* TG68K_FPU_ALU.vhd:1427:87  */
  assign n10528 = mant_result[0]; // extract
  /* TG68K_FPU_ALU.vhd:1427:97  */
  assign n10529 = n10528 | flags_inexact;
  /* TG68K_FPU_ALU.vhd:1427:73  */
  assign n10532 = n10529 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1427:73  */
  assign n10535 = n10529 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1420:65  */
  assign n10537 = operation_code == 7'b0100000;
  /* TG68K_FPU_ALU.vhd:1420:78  */
  assign n10539 = operation_code == 7'b0100100;
  /* TG68K_FPU_ALU.vhd:1420:78  */
  assign n10540 = n10537 | n10539;
  /* TG68K_FPU_ALU.vhd:1437:97  */
  assign n10541 = mant_result[0]; // extract
  /* TG68K_FPU_ALU.vhd:1439:73  */
  assign n10544 = flags_inexact ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1439:73  */
  assign n10547 = flags_inexact ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1434:65  */
  assign n10549 = operation_code == 7'b0000100;
  /* TG68K_FPU_ALU.vhd:1446:65  */
  assign n10551 = operation_code == 7'b0011000;
  /* TG68K_FPU_ALU.vhd:1446:78  */
  assign n10553 = operation_code == 7'b0011010;
  /* TG68K_FPU_ALU.vhd:1446:78  */
  assign n10554 = n10551 | n10553;
  /* TG68K_FPU_ALU.vhd:1446:88  */
  assign n10556 = operation_code == 7'b0000000;
  /* TG68K_FPU_ALU.vhd:1446:88  */
  assign n10557 = n10554 | n10556;
  /* TG68K_FPU_ALU.vhd:1454:92  */
  assign n10559 = $unsigned(exp_a) < $unsigned(15'b011111111111111);
  /* TG68K_FPU_ALU.vhd:1456:100  */
  assign n10560 = mant_a[63]; // extract
  /* TG68K_FPU_ALU.vhd:1457:100  */
  assign n10561 = mant_a[62]; // extract
  /* TG68K_FPU_ALU.vhd:1458:90  */
  assign n10562 = mant_a[61:0]; // extract
  /* TG68K_FPU_ALU.vhd:1458:104  */
  assign n10564 = n10562 != 62'b00000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1458:81  */
  assign n10567 = n10564 ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1454:73  */
  assign n10571 = n10559 ? n10560 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1454:73  */
  assign n10573 = n10559 ? n10561 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1454:73  */
  assign n10575 = n10559 ? n10567 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1451:65  */
  assign n10577 = operation_code == 7'b0000001;
  /* TG68K_FPU_ALU.vhd:1451:78  */
  assign n10579 = operation_code == 7'b0000011;
  /* TG68K_FPU_ALU.vhd:1451:78  */
  assign n10580 = n10577 | n10579;
  /* TG68K_FPU_ALU.vhd:1476:73  */
  assign n10583 = flags_inexact ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1476:73  */
  assign n10586 = flags_inexact ? 1'b1 : 1'b0;
  /* TG68K_FPU_ALU.vhd:1476:73  */
  assign n10589 = flags_inexact ? 1'b1 : 1'b0;
  assign n10590 = {n10580, n10557, n10549, n10540, n10526, n10516};
  /* TG68K_FPU_ALU.vhd:1396:57  */
  always @*
    case (n10590)
      6'b100000: n10592 = n10571;
      6'b010000: n10592 = 1'b0;
      6'b001000: n10592 = n10541;
      6'b000100: n10592 = n10527;
      6'b000010: n10592 = n10517;
      6'b000001: n10592 = n10509;
      default: n10592 = n10583;
    endcase
  /* TG68K_FPU_ALU.vhd:1396:57  */
  always @*
    case (n10590)
      6'b100000: n10594 = n10573;
      6'b010000: n10594 = 1'b0;
      6'b001000: n10594 = n10544;
      6'b000100: n10594 = n10532;
      6'b000010: n10594 = n10518;
      6'b000001: n10594 = n10511;
      default: n10594 = n10586;
    endcase
  /* TG68K_FPU_ALU.vhd:1396:57  */
  always @*
    case (n10590)
      6'b100000: n10597 = n10575;
      6'b010000: n10597 = 1'b0;
      6'b001000: n10597 = n10547;
      6'b000100: n10597 = n10535;
      6'b000010: n10597 = n10524;
      6'b000001: n10597 = 1'b0;
      default: n10597 = n10589;
    endcase
  /* TG68K_FPU_ALU.vhd:1493:113  */
  assign n10600 = round_bit | sticky_bit;
  /* TG68K_FPU_ALU.vhd:1493:147  */
  assign n10601 = mant_result[0]; // extract
  /* TG68K_FPU_ALU.vhd:1493:133  */
  assign n10602 = n10600 | n10601;
  /* TG68K_FPU_ALU.vhd:1493:92  */
  assign n10603 = n10602 & guard_bit;
  /* TG68K_FPU_ALU.vhd:1495:96  */
  assign n10605 = mant_result == 64'b1111111111111111111111111111111111111111111111111111111111111111;
  /* TG68K_FPU_ALU.vhd:1497:103  */
  assign n10607 = exp_result == 15'b111111111111110;
  /* TG68K_FPU_ALU.vhd:1503:122  */
  assign n10609 = exp_result + 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:1497:89  */
  assign n10611 = n10607 ? 15'b111111111111111 : n10609;
  /* TG68K_FPU_ALU.vhd:1497:89  */
  assign n10614 = n10607 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1493:73  */
  assign n10616 = n10624 ? 1'b1 : flags_overflow;
  /* TG68K_FPU_ALU.vhd:1507:116  */
  assign n10618 = mant_result + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1493:73  */
  assign n10619 = n10622 ? n10611 : n10501;
  /* TG68K_FPU_ALU.vhd:1495:81  */
  assign n10620 = n10605 ? n10614 : n10618;
  /* TG68K_FPU_ALU.vhd:1495:81  */
  assign n10621 = n10607 & n10605;
  /* TG68K_FPU_ALU.vhd:1493:73  */
  assign n10622 = n10605 & n10603;
  /* TG68K_FPU_ALU.vhd:1493:73  */
  assign n10623 = n10603 ? n10620 : n10502;
  /* TG68K_FPU_ALU.vhd:1493:73  */
  assign n10624 = n10621 & n10603;
  /* TG68K_FPU_ALU.vhd:1492:65  */
  assign n10626 = rounding_mode == 2'b00;
  /* TG68K_FPU_ALU.vhd:1510:65  */
  assign n10628 = rounding_mode == 2'b01;
  /* TG68K_FPU_ALU.vhd:1513:88  */
  assign n10629 = ~sign_result;
  /* TG68K_FPU_ALU.vhd:1513:115  */
  assign n10630 = guard_bit | round_bit;
  /* TG68K_FPU_ALU.vhd:1513:134  */
  assign n10631 = n10630 | sticky_bit;
  /* TG68K_FPU_ALU.vhd:1513:94  */
  assign n10632 = n10631 & n10629;
  /* TG68K_FPU_ALU.vhd:1515:96  */
  assign n10634 = mant_result == 64'b1111111111111111111111111111111111111111111111111111111111111111;
  /* TG68K_FPU_ALU.vhd:1516:103  */
  assign n10636 = exp_result == 15'b111111111111110;
  /* TG68K_FPU_ALU.vhd:1522:122  */
  assign n10638 = exp_result + 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:1516:89  */
  assign n10640 = n10636 ? 15'b111111111111111 : n10638;
  /* TG68K_FPU_ALU.vhd:1516:89  */
  assign n10643 = n10636 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1513:73  */
  assign n10645 = n10653 ? 1'b1 : flags_overflow;
  /* TG68K_FPU_ALU.vhd:1526:116  */
  assign n10647 = mant_result + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1513:73  */
  assign n10648 = n10651 ? n10640 : n10501;
  /* TG68K_FPU_ALU.vhd:1515:81  */
  assign n10649 = n10634 ? n10643 : n10647;
  /* TG68K_FPU_ALU.vhd:1515:81  */
  assign n10650 = n10636 & n10634;
  /* TG68K_FPU_ALU.vhd:1513:73  */
  assign n10651 = n10634 & n10632;
  /* TG68K_FPU_ALU.vhd:1513:73  */
  assign n10652 = n10632 ? n10649 : n10502;
  /* TG68K_FPU_ALU.vhd:1513:73  */
  assign n10653 = n10650 & n10632;
  /* TG68K_FPU_ALU.vhd:1512:65  */
  assign n10655 = rounding_mode == 2'b10;
  /* TG68K_FPU_ALU.vhd:1530:115  */
  assign n10656 = guard_bit | round_bit;
  /* TG68K_FPU_ALU.vhd:1530:134  */
  assign n10657 = n10656 | sticky_bit;
  /* TG68K_FPU_ALU.vhd:1530:94  */
  assign n10658 = n10657 & sign_result;
  /* TG68K_FPU_ALU.vhd:1532:96  */
  assign n10660 = mant_result == 64'b1111111111111111111111111111111111111111111111111111111111111111;
  /* TG68K_FPU_ALU.vhd:1533:103  */
  assign n10662 = exp_result == 15'b111111111111110;
  /* TG68K_FPU_ALU.vhd:1539:122  */
  assign n10664 = exp_result + 15'b000000000000001;
  /* TG68K_FPU_ALU.vhd:1533:89  */
  assign n10666 = n10662 ? 15'b111111111111111 : n10664;
  /* TG68K_FPU_ALU.vhd:1533:89  */
  assign n10669 = n10662 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b1000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU_ALU.vhd:1530:73  */
  assign n10671 = n10679 ? 1'b1 : flags_overflow;
  /* TG68K_FPU_ALU.vhd:1543:116  */
  assign n10673 = mant_result + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  /* TG68K_FPU_ALU.vhd:1530:73  */
  assign n10674 = n10677 ? n10666 : n10501;
  /* TG68K_FPU_ALU.vhd:1532:81  */
  assign n10675 = n10660 ? n10669 : n10673;
  /* TG68K_FPU_ALU.vhd:1532:81  */
  assign n10676 = n10662 & n10660;
  /* TG68K_FPU_ALU.vhd:1530:73  */
  assign n10677 = n10660 & n10658;
  /* TG68K_FPU_ALU.vhd:1530:73  */
  assign n10678 = n10658 ? n10675 : n10502;
  /* TG68K_FPU_ALU.vhd:1530:73  */
  assign n10679 = n10676 & n10658;
  /* TG68K_FPU_ALU.vhd:1529:65  */
  assign n10681 = rounding_mode == 2'b11;
  assign n10682 = {n10681, n10655, n10628, n10626};
  /* TG68K_FPU_ALU.vhd:1491:57  */
  always @*
    case (n10682)
      4'b1000: n10683 = n10674;
      4'b0100: n10683 = n10648;
      4'b0010: n10683 = n10501;
      4'b0001: n10683 = n10619;
      default: n10683 = n10501;
    endcase
  /* TG68K_FPU_ALU.vhd:1491:57  */
  always @*
    case (n10682)
      4'b1000: n10684 = n10678;
      4'b0100: n10684 = n10652;
      4'b0010: n10684 = n10502;
      4'b0001: n10684 = n10623;
      default: n10684 = n10502;
    endcase
  /* TG68K_FPU_ALU.vhd:1491:57  */
  always @*
    case (n10682)
      4'b1000: n10685 = n10671;
      4'b0100: n10685 = n10645;
      4'b0010: n10685 = flags_overflow;
      4'b0001: n10685 = n10616;
      default: n10685 = flags_overflow;
    endcase
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10686 = n9588 ? sign_result : n10493;
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10688 = n9588 ? 15'b000000000000000 : n10683;
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10690 = n9588 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n10684;
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10691 = n9588 ? guard_bit : n10592;
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10692 = n9588 ? round_bit : n10594;
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10693 = n9588 ? sticky_bit : n10597;
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10695 = n9588 ? flags_overflow : n10685;
  /* TG68K_FPU_ALU.vhd:1313:49  */
  assign n10697 = n9588 ? 1'b1 : n10503;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10699 = n9587 ? sign_result : n10686;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10701 = n9587 ? 15'b111111111111111 : n10688;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10703 = n9587 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n10690;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10704 = n9587 ? guard_bit : n10691;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10705 = n9587 ? round_bit : n10692;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10706 = n9587 ? sticky_bit : n10693;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10709 = n9587 ? 1'b1 : n10695;
  /* TG68K_FPU_ALU.vhd:1308:49  */
  assign n10710 = n9587 ? flags_underflow : n10697;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10712 = n9585 ? sign_result : n10699;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10714 = n9585 ? 15'b000000000000000 : n10701;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10716 = n9585 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n10703;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10717 = n9585 ? guard_bit : n10704;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10718 = n9585 ? round_bit : n10705;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10719 = n9585 ? sticky_bit : n10706;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10721 = n9585 ? flags_overflow : n10709;
  /* TG68K_FPU_ALU.vhd:1304:49  */
  assign n10722 = n9585 ? flags_underflow : n10710;
  /* TG68K_FPU_ALU.vhd:1301:41  */
  assign n10725 = alu_state == 3'b100;
  /* TG68K_FPU_ALU.vhd:1555:71  */
  assign n10726 = {sign_result, exp_result};
  /* TG68K_FPU_ALU.vhd:1555:84  */
  assign n10727 = {n10726, mant_result};
  /* TG68K_FPU_ALU.vhd:1553:41  */
  assign n10729 = alu_state == 3'b101;
  assign n10730 = {n10729, n10725, n9580, n7538, n7492, n7490};
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10732 = n10727;
      6'b010000: n10732 = n11054;
      6'b001000: n10732 = n11054;
      6'b000100: n10732 = n11054;
      6'b000010: n10732 = n11054;
      6'b000001: n10732 = n11054;
      default: n10732 = 80'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10736 = 1'b1;
      6'b010000: n10736 = n11056;
      6'b001000: n10736 = n11056;
      6'b000100: n10736 = n11056;
      6'b000010: n10736 = n11056;
      6'b000001: n10736 = 1'b0;
      default: n10736 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10739 = 1'b0;
      6'b010000: n10739 = n11058;
      6'b001000: n10739 = n11058;
      6'b000100: n10739 = n11058;
      6'b000010: n10739 = n11058;
      6'b000001: n10739 = n7485;
      default: n10739 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10743 = 1'b1;
      6'b010000: n10743 = n11060;
      6'b001000: n10743 = n11060;
      6'b000100: n10743 = n11060;
      6'b000010: n10743 = n11060;
      6'b000001: n10743 = 1'b0;
      default: n10743 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10745 = sign_a;
      6'b010000: n10745 = sign_a;
      6'b001000: n10745 = sign_a;
      6'b000100: n10745 = n7493;
      6'b000010: n10745 = sign_a;
      6'b000001: n10745 = sign_a;
      default: n10745 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10747 = sign_b;
      6'b010000: n10747 = sign_b;
      6'b001000: n10747 = sign_b;
      6'b000100: n10747 = n7496;
      6'b000010: n10747 = sign_b;
      6'b000001: n10747 = sign_b;
      default: n10747 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10749 = sign_result;
      6'b010000: n10749 = n10712;
      6'b001000: n10749 = n9555;
      6'b000100: n10749 = n7532;
      6'b000010: n10749 = sign_result;
      6'b000001: n10749 = sign_result;
      default: n10749 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10751 = exp_a;
      6'b010000: n10751 = exp_a;
      6'b001000: n10751 = exp_a;
      6'b000100: n10751 = n7494;
      6'b000010: n10751 = exp_a;
      6'b000001: n10751 = exp_a;
      default: n10751 = 15'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10753 = exp_b;
      6'b010000: n10753 = exp_b;
      6'b001000: n10753 = exp_b;
      6'b000100: n10753 = n7497;
      6'b000010: n10753 = exp_b;
      6'b000001: n10753 = exp_b;
      default: n10753 = 15'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10755 = exp_result;
      6'b010000: n10755 = n10714;
      6'b001000: n10755 = n9558;
      6'b000100: n10755 = n7533;
      6'b000010: n10755 = exp_result;
      6'b000001: n10755 = exp_result;
      default: n10755 = 15'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10757 = mant_a;
      6'b010000: n10757 = mant_a;
      6'b001000: n10757 = mant_a;
      6'b000100: n10757 = n7495;
      6'b000010: n10757 = mant_a;
      6'b000001: n10757 = mant_a;
      default: n10757 = 64'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10759 = mant_b;
      6'b010000: n10759 = mant_b;
      6'b001000: n10759 = mant_b;
      6'b000100: n10759 = n7498;
      6'b000010: n10759 = mant_b;
      6'b000001: n10759 = mant_b;
      default: n10759 = 64'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10761 = mant_result;
      6'b010000: n10761 = n10716;
      6'b001000: n10761 = n9561;
      6'b000100: n10761 = n7534;
      6'b000010: n10761 = mant_result;
      6'b000001: n10761 = mant_result;
      default: n10761 = 64'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10767 = 3'b000;
      6'b010000: n10767 = 3'b101;
      6'b001000: n10767 = 3'b100;
      6'b000100: n10767 = n7536;
      6'b000010: n10767 = 3'b010;
      6'b000001: n10767 = n7488;
      default: n10767 = 3'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10769 = mant_sum;
      6'b010000: n10769 = mant_sum;
      6'b001000: n10769 = n9562;
      6'b000100: n10769 = mant_sum;
      6'b000010: n10769 = mant_sum;
      6'b000001: n10769 = mant_sum;
      default: n10769 = 65'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10775 = mant_a_aligned;
      6'b010000: n10775 = mant_a_aligned;
      6'b001000: n10775 = n9565;
      6'b000100: n10775 = mant_a_aligned;
      6'b000010: n10775 = mant_a_aligned;
      6'b000001: n10775 = mant_a_aligned;
      default: n10775 = 65'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10777 = mant_b_aligned;
      6'b010000: n10777 = mant_b_aligned;
      6'b001000: n10777 = n9566;
      6'b000100: n10777 = mant_b_aligned;
      6'b000010: n10777 = mant_b_aligned;
      6'b000001: n10777 = mant_b_aligned;
      default: n10777 = 65'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10779 = exp_larger;
      6'b010000: n10779 = exp_larger;
      6'b001000: n10779 = n9567;
      6'b000100: n10779 = exp_larger;
      6'b000010: n10779 = exp_larger;
      6'b000001: n10779 = exp_larger;
      default: n10779 = 15'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10783 = guard_bit;
      6'b010000: n10783 = n10717;
      6'b001000: n10783 = guard_bit;
      6'b000100: n10783 = guard_bit;
      6'b000010: n10783 = guard_bit;
      6'b000001: n10783 = guard_bit;
      default: n10783 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10785 = round_bit;
      6'b010000: n10785 = n10718;
      6'b001000: n10785 = round_bit;
      6'b000100: n10785 = round_bit;
      6'b000010: n10785 = round_bit;
      6'b000001: n10785 = round_bit;
      default: n10785 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10787 = sticky_bit;
      6'b010000: n10787 = n10719;
      6'b001000: n10787 = sticky_bit;
      6'b000100: n10787 = sticky_bit;
      6'b000010: n10787 = sticky_bit;
      6'b000001: n10787 = sticky_bit;
      default: n10787 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10791 = mult_result;
      6'b010000: n10791 = mult_result;
      6'b001000: n10791 = n9569;
      6'b000100: n10791 = mult_result;
      6'b000010: n10791 = mult_result;
      6'b000001: n10791 = mult_result;
      default: n10791 = 128'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10793 = fmod_quotient;
      6'b010000: n10793 = fmod_quotient;
      6'b001000: n10793 = n9570;
      6'b000100: n10793 = fmod_quotient;
      6'b000010: n10793 = fmod_quotient;
      6'b000001: n10793 = fmod_quotient;
      default: n10793 = 8'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10796 = flags_overflow;
      6'b010000: n10796 = n10721;
      6'b001000: n10796 = n9571;
      6'b000100: n10796 = flags_overflow;
      6'b000010: n10796 = 1'b0;
      6'b000001: n10796 = flags_overflow;
      default: n10796 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10799 = flags_underflow;
      6'b010000: n10799 = n10722;
      6'b001000: n10799 = n9572;
      6'b000100: n10799 = flags_underflow;
      6'b000010: n10799 = 1'b0;
      6'b000001: n10799 = flags_underflow;
      default: n10799 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10802 = flags_inexact;
      6'b010000: n10802 = flags_inexact;
      6'b001000: n10802 = n9573;
      6'b000100: n10802 = flags_inexact;
      6'b000010: n10802 = 1'b0;
      6'b000001: n10802 = flags_inexact;
      default: n10802 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10805 = flags_invalid;
      6'b010000: n10805 = flags_invalid;
      6'b001000: n10805 = n9575;
      6'b000100: n10805 = flags_invalid;
      6'b000010: n10805 = 1'b0;
      6'b000001: n10805 = flags_invalid;
      default: n10805 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:283:33  */
  always @*
    case (n10730)
      6'b100000: n10808 = flags_div_by_zero;
      6'b010000: n10808 = flags_div_by_zero;
      6'b001000: n10808 = n9576;
      6'b000100: n10808 = flags_div_by_zero;
      6'b000010: n10808 = 1'b0;
      6'b000001: n10808 = flags_div_by_zero;
      default: n10808 = 1'bX;
    endcase
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10943 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10944 = clkena & n10943;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10945 = n10944 ? n10745 : sign_a;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10946 <= n10945;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10947 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10948 = clkena & n10947;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10949 = n10948 ? n10747 : sign_b;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10950 <= n10949;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10951 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10952 = clkena & n10951;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10953 = n10952 ? n10749 : sign_result;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10954 <= n10953;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10955 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10956 = clkena & n10955;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10957 = n10956 ? n10751 : exp_a;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10958 <= n10957;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10959 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10960 = clkena & n10959;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10961 = n10960 ? n10753 : exp_b;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10962 <= n10961;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10963 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10964 = clkena & n10963;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10965 = n10964 ? n10755 : exp_result;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10966 <= n10965;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10967 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10968 = clkena & n10967;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10969 = n10968 ? n10757 : mant_a;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10970 <= n10969;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10971 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10972 = clkena & n10971;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10973 = n10972 ? n10759 : mant_b;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10974 <= n10973;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10975 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10976 = clkena & n10975;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10977 = n10976 ? n10761 : mant_result;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10978 <= n10977;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10979 = clkena ? n10767 : alu_state;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n10980 <= 3'b000;
    else
      n10980 <= n10979;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10982 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10983 = clkena & n10982;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10984 = n10983 ? n10769 : mant_sum;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10985 <= n10984;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10995 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10996 = clkena & n10995;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n10997 = n10996 ? n10775 : mant_a_aligned;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n10998 <= n10997;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n10999 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11000 = clkena & n10999;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11001 = n11000 ? n10777 : mant_b_aligned;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n11002 <= n11001;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11003 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11004 = clkena & n11003;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11005 = n11004 ? n10779 : exp_larger;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n11006 <= n11005;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11011 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11012 = clkena & n11011;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11013 = n11012 ? n10783 : guard_bit;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n11014 <= n11013;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11015 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11016 = clkena & n11015;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11017 = n11016 ? n10785 : round_bit;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n11018 <= n11017;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11019 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11020 = clkena & n11019;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11021 = n11020 ? n10787 : sticky_bit;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n11022 <= n11021;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11029 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11030 = clkena & n11029;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11031 = n11030 ? n10791 : mult_result;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n11032 <= n11031;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11039 = ~n7481;
  /* TG68K_FPU_ALU.vhd:262:9  */
  assign n11040 = clkena & n11039;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11041 = n11040 ? n10793 : fmod_quotient;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk)
    n11042 <= n11041;
  initial
    n11042 = 8'b00000000;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11043 = clkena ? n10796 : flags_overflow;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11044 <= 1'b0;
    else
      n11044 <= n11043;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11045 = clkena ? n10799 : flags_underflow;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11046 <= 1'b0;
    else
      n11046 <= n11045;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11047 = clkena ? n10802 : flags_inexact;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11048 <= 1'b0;
    else
      n11048 <= n11047;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11049 = clkena ? n10805 : flags_invalid;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11050 <= 1'b0;
    else
      n11050 <= n11049;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11051 = clkena ? n10808 : flags_div_by_zero;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11052 <= 1'b0;
    else
      n11052 <= n11051;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11053 = clkena ? n10732 : n11054;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11054 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n11054 <= n11053;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11055 = clkena ? n10736 : n11056;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11056 <= 1'b0;
    else
      n11056 <= n11055;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11057 = clkena ? n10739 : n11058;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11058 <= 1'b0;
    else
      n11058 <= n11057;
  /* TG68K_FPU_ALU.vhd:281:17  */
  assign n11059 = clkena ? n10743 : n11060;
  /* TG68K_FPU_ALU.vhd:281:17  */
  always @(posedge clk or posedge n7481)
    if (n7481)
      n11060 <= 1'b0;
    else
      n11060 <= n11059;
endmodule

module tg68k_fpu_decoder
  (input  clk,
   input  nreset,
   input  [15:0] opcode,
   input  [15:0] extension_word,
   input  decode_enable,
   output [3:0] instruction_type,
   output [6:0] operation_code,
   output [2:0] source_format,
   output [2:0] dest_format,
   output [2:0] source_reg,
   output [2:0] dest_reg,
   output [2:0] ea_mode,
   output [2:0] ea_register,
   output needs_extension_word,
   output valid_instruction,
   output privileged_instruction,
   output illegal_instruction,
   output unsupported_instruction);
  wire [2:0] coprocessor_id;
  wire [2:0] inst_type_bits;
  wire [2:0] format_field;
  wire [6:0] opmode_field;
  wire [2:0] rm_field;
  wire [2:0] rn_field;
  wire [3:0] instruction_type_int;
  wire valid_f_line;
  wire valid_coprocessor_id;
  wire valid_format;
  wire valid_opmode;
  wire [2:0] n7117;
  wire [2:0] n7118;
  wire [2:0] n7119;
  wire [2:0] n7120;
  wire n7122;
  wire [2:0] n7123;
  wire [6:0] n7124;
  wire [2:0] n7125;
  wire [2:0] n7126;
  wire [2:0] n7128;
  wire [6:0] n7130;
  wire [2:0] n7132;
  wire [2:0] n7134;
  wire [3:0] n7137;
  wire n7139;
  wire n7141;
  wire n7142;
  wire [2:0] n7143;
  wire n7145;
  wire [2:0] n7146;
  wire n7148;
  wire n7149;
  wire [2:0] n7150;
  wire n7152;
  wire [2:0] n7153;
  wire n7155;
  wire n7156;
  wire n7157;
  wire [3:0] n7160;
  wire n7162;
  wire [2:0] n7163;
  wire n7165;
  wire [2:0] n7166;
  wire n7168;
  wire [2:0] n7169;
  wire n7171;
  wire [2:0] n7172;
  wire n7174;
  wire n7175;
  wire [3:0] n7178;
  wire [3:0] n7180;
  wire [3:0] n7182;
  wire n7184;
  wire n7186;
  wire n7188;
  wire n7190;
  wire n7192;
  wire n7193;
  wire n7194;
  wire [7:0] n7195;
  wire n7197;
  wire n7198;
  wire n7199;
  wire n7200;
  wire n7201;
  wire [2:0] n7202;
  wire n7204;
  wire [7:0] n7205;
  wire n7207;
  wire n7208;
  wire [4:0] n7209;
  wire n7211;
  wire [3:0] n7214;
  wire n7217;
  wire [3:0] n7219;
  wire n7221;
  wire [3:0] n7223;
  wire n7225;
  wire [3:0] n7227;
  wire n7229;
  wire [2:0] n7230;
  wire n7232;
  wire n7235;
  wire [3:0] n7238;
  wire n7240;
  wire [7:0] n7241;
  reg n7251;
  reg n7255;
  reg [3:0] n7261;
  wire n7263;
  wire n7266;
  wire [3:0] n7269;
  wire [3:0] n7273;
  wire n7275;
  wire n7278;
  wire n7280;
  wire n7283;
  wire n7285;
  wire n7287;
  wire n7288;
  wire n7290;
  wire n7291;
  wire n7293;
  wire n7294;
  wire n7296;
  wire n7297;
  wire n7299;
  wire n7300;
  wire n7302;
  wire n7303;
  reg n7306;
  wire n7308;
  wire n7310;
  wire n7311;
  wire n7313;
  wire n7315;
  wire n7316;
  wire n7317;
  wire n7319;
  wire n7321;
  wire n7322;
  wire n7323;
  wire n7326;
  wire n7327;
  wire n7328;
  wire n7329;
  wire n7330;
  wire n7331;
  wire n7332;
  wire n7333;
  wire n7334;
  wire n7335;
  localparam n7337 = 1'b0;
  wire n7339;
  wire [2:0] n7340;
  localparam [2:0] n7342 = 3'b010;
  assign instruction_type = instruction_type_int; //(module output)
  assign operation_code = opmode_field; //(module output)
  assign source_format = n7340; //(module output)
  assign dest_format = n7342; //(module output)
  assign source_reg = rm_field; //(module output)
  assign dest_reg = rn_field; //(module output)
  assign ea_mode = n7119; //(module output)
  assign ea_register = n7120; //(module output)
  assign needs_extension_word = n7263; //(module output)
  assign valid_instruction = n7330; //(module output)
  assign privileged_instruction = n7266; //(module output)
  assign illegal_instruction = n7335; //(module output)
  assign unsupported_instruction = n7337; //(module output)
  /* TG68K_FPU_Decoder.vhd:85:16  */
  assign coprocessor_id = n7117; // (signal)
  /* TG68K_FPU_Decoder.vhd:86:16  */
  assign inst_type_bits = n7118; // (signal)
  /* TG68K_FPU_Decoder.vhd:87:16  */
  assign format_field = n7128; // (signal)
  /* TG68K_FPU_Decoder.vhd:88:16  */
  assign opmode_field = n7130; // (signal)
  /* TG68K_FPU_Decoder.vhd:89:16  */
  assign rm_field = n7132; // (signal)
  /* TG68K_FPU_Decoder.vhd:90:16  */
  assign rn_field = n7134; // (signal)
  /* TG68K_FPU_Decoder.vhd:91:16  */
  assign instruction_type_int = n7269; // (signal)
  /* TG68K_FPU_Decoder.vhd:94:16  */
  assign valid_f_line = n7278; // (signal)
  /* TG68K_FPU_Decoder.vhd:95:16  */
  assign valid_coprocessor_id = n7283; // (signal)
  /* TG68K_FPU_Decoder.vhd:96:16  */
  assign valid_format = n7306; // (signal)
  /* TG68K_FPU_Decoder.vhd:97:16  */
  assign valid_opmode = n7326; // (signal)
  /* TG68K_FPU_Decoder.vhd:110:41  */
  assign n7117 = opcode[11:9]; // extract
  /* TG68K_FPU_Decoder.vhd:111:41  */
  assign n7118 = opcode[8:6]; // extract
  /* TG68K_FPU_Decoder.vhd:112:34  */
  assign n7119 = opcode[5:3]; // extract
  /* TG68K_FPU_Decoder.vhd:113:38  */
  assign n7120 = opcode[2:0]; // extract
  /* TG68K_FPU_Decoder.vhd:124:35  */
  assign n7122 = inst_type_bits == 3'b000;
  /* TG68K_FPU_Decoder.vhd:127:55  */
  assign n7123 = extension_word[12:10]; // extract
  /* TG68K_FPU_Decoder.vhd:128:55  */
  assign n7124 = extension_word[6:0]; // extract
  /* TG68K_FPU_Decoder.vhd:129:51  */
  assign n7125 = extension_word[15:13]; // extract
  /* TG68K_FPU_Decoder.vhd:130:51  */
  assign n7126 = extension_word[2:0]; // extract
  /* TG68K_FPU_Decoder.vhd:124:17  */
  assign n7128 = n7122 ? n7123 : 3'b000;
  /* TG68K_FPU_Decoder.vhd:124:17  */
  assign n7130 = n7122 ? n7124 : 7'b0000000;
  /* TG68K_FPU_Decoder.vhd:124:17  */
  assign n7132 = n7122 ? n7125 : 3'b000;
  /* TG68K_FPU_Decoder.vhd:124:17  */
  assign n7134 = n7122 ? n7126 : 3'b000;
  /* TG68K_FPU_Decoder.vhd:147:26  */
  assign n7137 = opcode[15:12]; // extract
  /* TG68K_FPU_Decoder.vhd:147:41  */
  assign n7139 = n7137 == 4'b1111;
  /* TG68K_FPU_Decoder.vhd:147:69  */
  assign n7141 = coprocessor_id == 3'b001;
  /* TG68K_FPU_Decoder.vhd:147:50  */
  assign n7142 = n7141 & n7139;
  /* TG68K_FPU_Decoder.vhd:153:51  */
  assign n7143 = opcode[5:3]; // extract
  /* TG68K_FPU_Decoder.vhd:153:64  */
  assign n7145 = n7143 == 3'b010;
  /* TG68K_FPU_Decoder.vhd:153:82  */
  assign n7146 = opcode[2:0]; // extract
  /* TG68K_FPU_Decoder.vhd:153:95  */
  assign n7148 = n7146 == 3'b101;
  /* TG68K_FPU_Decoder.vhd:153:72  */
  assign n7149 = n7148 & n7145;
  /* TG68K_FPU_Decoder.vhd:154:51  */
  assign n7150 = opcode[5:3]; // extract
  /* TG68K_FPU_Decoder.vhd:154:64  */
  assign n7152 = n7150 == 3'b001;
  /* TG68K_FPU_Decoder.vhd:154:82  */
  assign n7153 = opcode[2:0]; // extract
  /* TG68K_FPU_Decoder.vhd:154:95  */
  assign n7155 = n7153 == 3'b101;
  /* TG68K_FPU_Decoder.vhd:154:72  */
  assign n7156 = n7155 & n7152;
  /* TG68K_FPU_Decoder.vhd:153:104  */
  assign n7157 = n7149 | n7156;
  /* TG68K_FPU_Decoder.vhd:153:41  */
  assign n7160 = n7157 ? 4'b0011 : 4'b0000;
  /* TG68K_FPU_Decoder.vhd:149:33  */
  assign n7162 = inst_type_bits == 3'b000;
  /* TG68K_FPU_Decoder.vhd:167:50  */
  assign n7163 = opcode[5:3]; // extract
  /* TG68K_FPU_Decoder.vhd:167:63  */
  assign n7165 = n7163 == 3'b001;
  /* TG68K_FPU_Decoder.vhd:169:53  */
  assign n7166 = opcode[5:3]; // extract
  /* TG68K_FPU_Decoder.vhd:169:66  */
  assign n7168 = n7166 == 3'b111;
  /* TG68K_FPU_Decoder.vhd:170:58  */
  assign n7169 = opcode[2:0]; // extract
  /* TG68K_FPU_Decoder.vhd:170:71  */
  assign n7171 = n7169 == 3'b010;
  /* TG68K_FPU_Decoder.vhd:170:88  */
  assign n7172 = opcode[2:0]; // extract
  /* TG68K_FPU_Decoder.vhd:170:101  */
  assign n7174 = n7172 == 3'b011;
  /* TG68K_FPU_Decoder.vhd:170:79  */
  assign n7175 = n7171 | n7174;
  /* TG68K_FPU_Decoder.vhd:170:49  */
  assign n7178 = n7175 ? 4'b1000 : 4'b0101;
  /* TG68K_FPU_Decoder.vhd:169:41  */
  assign n7180 = n7168 ? n7178 : 4'b0101;
  /* TG68K_FPU_Decoder.vhd:167:41  */
  assign n7182 = n7165 ? 4'b0101 : n7180;
  /* TG68K_FPU_Decoder.vhd:166:33  */
  assign n7184 = inst_type_bits == 3'b001;
  /* TG68K_FPU_Decoder.vhd:180:33  */
  assign n7186 = inst_type_bits == 3'b010;
  /* TG68K_FPU_Decoder.vhd:184:33  */
  assign n7188 = inst_type_bits == 3'b011;
  /* TG68K_FPU_Decoder.vhd:188:33  */
  assign n7190 = inst_type_bits == 3'b100;
  /* TG68K_FPU_Decoder.vhd:193:33  */
  assign n7192 = inst_type_bits == 3'b101;
  /* TG68K_FPU_Decoder.vhd:199:58  */
  assign n7193 = extension_word[15]; // extract
  /* TG68K_FPU_Decoder.vhd:199:63  */
  assign n7194 = ~n7193;
  /* TG68K_FPU_Decoder.vhd:203:59  */
  assign n7195 = opcode[15:8]; // extract
  /* TG68K_FPU_Decoder.vhd:203:73  */
  assign n7197 = n7195 == 8'b11110010;
  /* TG68K_FPU_Decoder.vhd:204:67  */
  assign n7198 = extension_word[15]; // extract
  /* TG68K_FPU_Decoder.vhd:203:82  */
  assign n7199 = n7198 & n7197;
  /* TG68K_FPU_Decoder.vhd:205:67  */
  assign n7200 = extension_word[14]; // extract
  /* TG68K_FPU_Decoder.vhd:204:79  */
  assign n7201 = n7200 & n7199;
  /* TG68K_FPU_Decoder.vhd:207:74  */
  assign n7202 = extension_word[12:10]; // extract
  /* TG68K_FPU_Decoder.vhd:207:89  */
  assign n7204 = n7202 != 3'b000;
  /* TG68K_FPU_Decoder.vhd:207:116  */
  assign n7205 = extension_word[7:0]; // extract
  /* TG68K_FPU_Decoder.vhd:207:129  */
  assign n7207 = n7205 == 8'b00000000;
  /* TG68K_FPU_Decoder.vhd:207:98  */
  assign n7208 = n7207 & n7204;
  /* TG68K_FPU_Decoder.vhd:210:77  */
  assign n7209 = extension_word[12:8]; // extract
  /* TG68K_FPU_Decoder.vhd:210:91  */
  assign n7211 = n7209 == 5'b00000;
  /* TG68K_FPU_Decoder.vhd:210:57  */
  assign n7214 = n7211 ? 4'b0011 : 4'b0000;
  /* TG68K_FPU_Decoder.vhd:207:57  */
  assign n7217 = n7208 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:207:57  */
  assign n7219 = n7208 ? 4'b1001 : n7214;
  /* TG68K_FPU_Decoder.vhd:203:49  */
  assign n7221 = n7201 ? n7217 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:203:49  */
  assign n7223 = n7201 ? n7219 : 4'b0000;
  /* TG68K_FPU_Decoder.vhd:199:41  */
  assign n7225 = n7194 ? 1'b0 : n7221;
  /* TG68K_FPU_Decoder.vhd:199:41  */
  assign n7227 = n7194 ? 4'b0001 : n7223;
  /* TG68K_FPU_Decoder.vhd:198:33  */
  assign n7229 = inst_type_bits == 3'b110;
  /* TG68K_FPU_Decoder.vhd:224:58  */
  assign n7230 = extension_word[15:13]; // extract
  /* TG68K_FPU_Decoder.vhd:224:73  */
  assign n7232 = n7230 == 3'b100;
  /* TG68K_FPU_Decoder.vhd:224:41  */
  assign n7235 = n7232 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:224:41  */
  assign n7238 = n7232 ? 4'b0100 : 4'b0010;
  /* TG68K_FPU_Decoder.vhd:223:33  */
  assign n7240 = inst_type_bits == 3'b111;
  assign n7241 = {n7240, n7229, n7192, n7190, n7188, n7186, n7184, n7162};
  /* TG68K_FPU_Decoder.vhd:148:25  */
  always @*
    case (n7241)
      8'b10000000: n7251 = 1'b1;
      8'b01000000: n7251 = 1'b1;
      8'b00100000: n7251 = 1'b0;
      8'b00010000: n7251 = 1'b0;
      8'b00001000: n7251 = 1'b1;
      8'b00000100: n7251 = 1'b1;
      8'b00000010: n7251 = 1'b1;
      8'b00000001: n7251 = 1'b1;
      default: n7251 = 1'b1;
    endcase
  /* TG68K_FPU_Decoder.vhd:148:25  */
  always @*
    case (n7241)
      8'b10000000: n7255 = n7235;
      8'b01000000: n7255 = n7225;
      8'b00100000: n7255 = 1'b1;
      8'b00010000: n7255 = 1'b1;
      8'b00001000: n7255 = 1'b0;
      8'b00000100: n7255 = 1'b0;
      8'b00000010: n7255 = 1'b0;
      8'b00000001: n7255 = 1'b0;
      default: n7255 = 1'b0;
    endcase
  /* TG68K_FPU_Decoder.vhd:148:25  */
  always @*
    case (n7241)
      8'b10000000: n7261 = n7238;
      8'b01000000: n7261 = n7227;
      8'b00100000: n7261 = 4'b0111;
      8'b00010000: n7261 = 4'b0110;
      8'b00001000: n7261 = 4'b0101;
      8'b00000100: n7261 = 4'b0101;
      8'b00000010: n7261 = n7182;
      8'b00000001: n7261 = n7160;
      default: n7261 = 4'b0000;
    endcase
  /* TG68K_FPU_Decoder.vhd:147:17  */
  assign n7263 = n7142 ? n7251 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:147:17  */
  assign n7266 = n7142 ? n7255 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:147:17  */
  assign n7269 = n7142 ? n7261 : 4'b0000;
  /* TG68K_FPU_Decoder.vhd:246:26  */
  assign n7273 = opcode[15:12]; // extract
  /* TG68K_FPU_Decoder.vhd:246:41  */
  assign n7275 = n7273 == 4'b1111;
  /* TG68K_FPU_Decoder.vhd:246:17  */
  assign n7278 = n7275 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:253:35  */
  assign n7280 = coprocessor_id == 3'b001;
  /* TG68K_FPU_Decoder.vhd:253:17  */
  assign n7283 = n7280 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:261:25  */
  assign n7285 = format_field == 3'b000;
  /* TG68K_FPU_Decoder.vhd:261:42  */
  assign n7287 = format_field == 3'b001;
  /* TG68K_FPU_Decoder.vhd:261:42  */
  assign n7288 = n7285 | n7287;
  /* TG68K_FPU_Decoder.vhd:261:58  */
  assign n7290 = format_field == 3'b010;
  /* TG68K_FPU_Decoder.vhd:261:58  */
  assign n7291 = n7288 | n7290;
  /* TG68K_FPU_Decoder.vhd:261:76  */
  assign n7293 = format_field == 3'b011;
  /* TG68K_FPU_Decoder.vhd:261:76  */
  assign n7294 = n7291 | n7293;
  /* TG68K_FPU_Decoder.vhd:262:48  */
  assign n7296 = format_field == 3'b100;
  /* TG68K_FPU_Decoder.vhd:262:48  */
  assign n7297 = n7294 | n7296;
  /* TG68K_FPU_Decoder.vhd:262:62  */
  assign n7299 = format_field == 3'b101;
  /* TG68K_FPU_Decoder.vhd:262:62  */
  assign n7300 = n7297 | n7299;
  /* TG68K_FPU_Decoder.vhd:262:78  */
  assign n7302 = format_field == 3'b110;
  /* TG68K_FPU_Decoder.vhd:262:78  */
  assign n7303 = n7300 | n7302;
  /* TG68K_FPU_Decoder.vhd:260:17  */
  always @*
    case (n7303)
      1'b1: n7306 = 1'b1;
      default: n7306 = 1'b0;
    endcase
  /* TG68K_FPU_Decoder.vhd:271:34  */
  assign n7308 = $unsigned(opmode_field) >= $unsigned(7'b0000000);
  /* TG68K_FPU_Decoder.vhd:271:64  */
  assign n7310 = $unsigned(opmode_field) <= $unsigned(7'b0001111);
  /* TG68K_FPU_Decoder.vhd:271:47  */
  assign n7311 = n7310 & n7308;
  /* TG68K_FPU_Decoder.vhd:272:34  */
  assign n7313 = $unsigned(opmode_field) >= $unsigned(7'b0100000);
  /* TG68K_FPU_Decoder.vhd:272:64  */
  assign n7315 = $unsigned(opmode_field) <= $unsigned(7'b0101111);
  /* TG68K_FPU_Decoder.vhd:272:47  */
  assign n7316 = n7315 & n7313;
  /* TG68K_FPU_Decoder.vhd:271:78  */
  assign n7317 = n7311 | n7316;
  /* TG68K_FPU_Decoder.vhd:273:34  */
  assign n7319 = $unsigned(opmode_field) >= $unsigned(7'b0001100);
  /* TG68K_FPU_Decoder.vhd:273:64  */
  assign n7321 = $unsigned(opmode_field) <= $unsigned(7'b0011111);
  /* TG68K_FPU_Decoder.vhd:273:47  */
  assign n7322 = n7321 & n7319;
  /* TG68K_FPU_Decoder.vhd:272:78  */
  assign n7323 = n7317 | n7322;
  /* TG68K_FPU_Decoder.vhd:271:17  */
  assign n7326 = n7323 ? 1'b1 : 1'b0;
  /* TG68K_FPU_Decoder.vhd:280:52  */
  assign n7327 = decode_enable & valid_f_line;
  /* TG68K_FPU_Decoder.vhd:280:69  */
  assign n7328 = n7327 & valid_coprocessor_id;
  /* TG68K_FPU_Decoder.vhd:280:94  */
  assign n7329 = n7328 & valid_format;
  /* TG68K_FPU_Decoder.vhd:280:111  */
  assign n7330 = n7329 & valid_opmode;
  /* TG68K_FPU_Decoder.vhd:281:76  */
  assign n7331 = valid_f_line & valid_coprocessor_id;
  /* TG68K_FPU_Decoder.vhd:281:101  */
  assign n7332 = n7331 & valid_format;
  /* TG68K_FPU_Decoder.vhd:281:118  */
  assign n7333 = n7332 & valid_opmode;
  /* TG68K_FPU_Decoder.vhd:281:58  */
  assign n7334 = ~n7333;
  /* TG68K_FPU_Decoder.vhd:281:54  */
  assign n7335 = decode_enable & n7334;
  /* TG68K_FPU_Decoder.vhd:294:65  */
  assign n7339 = instruction_type_int == 4'b0000;
  /* TG68K_FPU_Decoder.vhd:294:39  */
  assign n7340 = n7339 ? format_field : 3'b010;
endmodule

module TG68K_FPU
  (input  clk,
   input  nReset,
   input  clkena,
   input  [15:0] opcode,
   input  [15:0] extension_word,
   input  fpu_enable,
   input  supervisor_mode,
   input  [31:0] cpu_data_in,
   input  [31:0] cpu_address_in,
   input  fsave_data_request,
   input  [5:0] fsave_data_index,
   input  frestore_data_write,
   input  [31:0] frestore_data_in,
   input  fmovem_data_request,
   input  [2:0] fmovem_reg_index,
   input  fmovem_data_write,
   input  [79:0] fmovem_data_in,
   input  [4:0] cir_address,
   input  cir_write,
   input  cir_read,
   input  [15:0] cir_data_in,
   output [31:0] fpu_data_out,
   output [79:0] fmovem_data_out,
   output fpu_busy,
   output fpu_done,
   output fpu_exception,
   output [7:0] exception_code,
   output [31:0] fpcr_out,
   output [31:0] fpsr_out,
   output [31:0] fpiar_out,
   output [7:0] fsave_frame_size,
   output fsave_size_valid,
   output [15:0] cir_data_out,
   output cir_data_valid);
  reg fpu_done_i;
  reg fpu_exception_i;
  reg cir_data_valid_i;
  wire [639:0] fp_registers;
  reg fp_reg_write_enable;
  reg [2:0] fp_reg_write_addr;
  reg [79:0] fp_reg_write_data;
  reg fp_reg_access_valid;
  reg [31:0] fpcr;
  reg [31:0] fpsr;
  reg [31:0] fpiar;
  reg fpcr_rounding_mode_valid;
  reg fpcr_precision_valid;
  wire [1:0] fpcr_precision_bits;
  reg [15:0] response_cir;
  reg [15:0] command_cir;
  reg [15:0] condition_cir;
  reg [15:0] save_cir;
  reg cir_read_reg;
  reg cir_write_reg;
  reg cir_read_active;
  reg [9:0] cir_timeout_counter;
  reg [9:0] state_timeout_counter;
  reg command_pending;
  reg command_valid;
  reg restore_privilege_violation;
  reg cir_address_error;
  reg [2:0] current_privilege_level;
  reg [2:0] cir_handshake_state;
  reg [15:0] operation_word_cir;
  reg [31:0] command_address_cir;
  reg [3:0] fpu_state;
  reg fpu_busy_internal;
  wire [7:0] fsave_frame_format;
  reg [7:0] fsave_frame_size_internal;
  reg fsave_size_valid_internal;
  reg [7:0] fsave_frame_format_latched;
  reg fpu_just_reset;
  wire [7:0] movem_register_list;
  wire movem_direction;
  reg [7:0] timeout_counter;
  reg [5:0] fsave_counter;
  wire [7:0] frestore_frame_format;
  wire [639:0] frestore_fp_temp;
  wire [3:0] decoder_instruction_type;
  wire [6:0] decoder_operation_code;
  wire [2:0] decoder_source_format;
  wire [2:0] decoder_dest_format;
  wire [2:0] decoder_source_reg;
  wire [2:0] decoder_dest_reg;
  wire [2:0] decoder_ea_mode;
  wire [2:0] decoder_ea_register;
  wire decoder_valid_instruction;
  wire decoder_illegal;
  wire decoder_unsupported;
  wire [6:0] fpu_operation;
  wire [2:0] source_reg;
  wire [2:0] dest_reg;
  wire [2:0] data_format;
  wire [2:0] ea_mode;
  wire [2:0] ea_register;
  wire [7:0] exception_code_internal;
  wire alu_start_operation;
  wire [6:0] alu_operation_code;
  wire [79:0] alu_operand_a;
  wire [79:0] alu_operand_b;
  wire [79:0] alu_result;
  wire alu_result_valid;
  wire alu_overflow;
  wire alu_underflow;
  wire alu_inexact;
  wire exception_reset;
  wire exception_op_valid;
  wire [7:0] exception_op_type;
  wire alu_invalid;
  wire alu_divide_by_zero;
  wire alu_operation_done;
  wire [7:0] alu_quotient_byte;
  wire trans_start_operation;
  wire [6:0] trans_operation_code;
  wire [79:0] trans_operand;
  wire [79:0] trans_result;
  wire trans_result_valid;
  wire trans_overflow;
  wire trans_underflow;
  wire trans_inexact;
  wire trans_invalid;
  wire trans_operation_done;
  wire [79:0] final_result;
  wire final_overflow;
  wire final_underflow;
  wire final_inexact;
  wire final_invalid;
  wire [79:0] result_data;
  wire converter_start;
  wire [2:0] converter_source_format;
  wire [2:0] converter_dest_format;
  wire [95:0] converter_data_in;
  wire [6:0] rom_offset;
  wire rom_read_enable;
  wire [79:0] constrom_result;
  wire constrom_valid;
  wire movem_start;
  wire movem_done;
  reg movem_predecrement;
  reg movem_postincrement;
  wire [2:0] movem_reg_address;
  wire [79:0] movem_reg_data_in;
  wire movem_unit_address_error;
  wire [5:0] fp_to_int_shift;
  wire [31:0] fp_to_int_result;
  wire [31:0] exception_fpsr_out;
  wire exception_pending_internal;
  wire [7:0] exception_vector_internal;
  wire [79:0] exception_corrected_result;
  wire [3:0] fpu_decoder_n81;
  wire [6:0] fpu_decoder_n82;
  wire [2:0] fpu_decoder_n83;
  wire [2:0] fpu_decoder_n84;
  wire [2:0] fpu_decoder_n85;
  wire [2:0] fpu_decoder_n86;
  wire [2:0] fpu_decoder_n87;
  wire [2:0] fpu_decoder_n88;
  wire fpu_decoder_n90;
  wire fpu_decoder_n92;
  wire fpu_decoder_n93;
  wire \fpu_decoder.needs_extension_word ;
  wire \fpu_decoder.privileged_instruction ;
  wire \fpu_alu.operation_busy ;
  wire [1:0] n118;
  wire [79:0] fpu_trans_n129;
  wire fpu_trans_n130;
  wire fpu_trans_n131;
  wire fpu_trans_n132;
  wire fpu_trans_n133;
  wire fpu_trans_n134;
  wire fpu_trans_n136;
  wire \fpu_trans.operation_busy ;
  wire \fpu_converter.conversion_done ;
  wire \fpu_converter.conversion_valid ;
  wire [79:0] \fpu_converter.data_out ;
  wire \fpu_converter.overflow ;
  wire \fpu_converter.underflow ;
  wire \fpu_converter.inexact ;
  wire \fpu_converter.invalid ;
  wire [79:0] fpu_const_rom_n173;
  wire fpu_const_rom_n174;
  wire \fpu_movem.movem_busy ;
  wire [79:0] \fpu_movem.fmovem_data_out ;
  wire [79:0] \fpu_movem.reg_data_out ;
  wire \fpu_movem.reg_write_enable ;
  wire n190;
  wire n191;
  wire [7:0] n193;
  wire n194;
  wire n195;
  wire [31:0] n196;
  wire [7:0] n197;
  wire [79:0] n202;
  wire n204;
  wire n207;
  wire [79:0] n209;
  wire n211;
  wire n213;
  wire [79:0] n214;
  wire n216;
  wire n218;
  wire [79:0] n219;
  wire n221;
  wire n223;
  wire [79:0] n224;
  wire n226;
  wire n228;
  wire [79:0] n229;
  wire n231;
  wire n233;
  wire [79:0] n234;
  wire n236;
  wire n238;
  wire [79:0] n239;
  wire n241;
  wire n243;
  wire n245;
  wire n247;
  wire n248;
  wire n251;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n271;
  wire n272;
  wire n273;
  wire [7:0] n276;
  wire [7:0] n279;
  wire [7:0] n281;
  wire [7:0] n283;
  wire [7:0] n285;
  wire [7:0] n287;
  wire n294;
  wire [6:0] n297;
  wire [2:0] n299;
  wire [2:0] n301;
  wire [2:0] n303;
  wire [2:0] n305;
  wire [2:0] n307;
  wire n743;
  wire n745;
  wire [30:0] n746;
  wire [31:0] n747;
  wire n749;
  wire [2:0] n752;
  wire [639:0] n755;
  wire n756;
  wire n757;
  wire [31:0] n759;
  wire [31:0] n761;
  wire n763;
  wire n766;
  wire [3:0] n769;
  wire [7:0] n771;
  wire [5:0] n773;
  wire [7:0] n775;
  wire n776;
  wire n778;
  wire n781;
  wire [3:0] n784;
  wire [5:0] n786;
  wire [7:0] n788;
  wire [7:0] n794;
  wire n795;
  wire n797;
  wire n799;
  wire n801;
  wire [2:0] n802;
  reg n805;
  reg n808;
  reg [3:0] n812;
  wire n813;
  wire n814;
  wire n817;
  wire [3:0] n819;
  wire [7:0] n821;
  wire n822;
  wire n823;
  wire [3:0] n824;
  wire [7:0] n825;
  wire n826;
  wire n828;
  wire [3:0] n830;
  wire [7:0] n831;
  wire n832;
  wire n833;
  wire [3:0] n834;
  wire [5:0] n835;
  wire [7:0] n836;
  wire [7:0] n839;
  wire [31:0] n841;
  wire n843;
  wire n844;
  wire [3:0] n846;
  wire [7:0] n848;
  wire [5:0] n849;
  wire [7:0] n850;
  wire [7:0] n853;
  wire n855;
  wire n857;
  wire n859;
  wire [3:0] n861;
  wire [7:0] n863;
  wire n865;
  wire n867;
  wire n868;
  wire n870;
  wire n871;
  wire n873;
  wire n875;
  wire [3:0] n877;
  wire [7:0] n879;
  wire n881;
  wire n883;
  wire n884;
  reg n885;
  reg n886;
  reg [3:0] n887;
  reg [7:0] n888;
  wire n890;
  wire n892;
  wire n894;
  wire n896;
  wire [3:0] n898;
  wire [7:0] n900;
  wire n902;
  wire n904;
  wire [3:0] n906;
  wire [7:0] n908;
  wire [2:0] n909;
  reg n910;
  reg n911;
  reg [3:0] n912;
  reg [7:0] n913;
  wire n915;
  wire n917;
  wire n918;
  wire [31:0] n919;
  wire n920;
  wire n922;
  wire n935;
  wire n937;
  wire n941;
  wire [4:0] n943;
  wire n945;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n972;
  wire n973;
  wire n975;
  wire n977;
  wire n978;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n995;
  wire n996;
  wire n997;
  wire n999;
  wire n1000;
  wire n1002;
  wire n1004;
  wire [15:0] n1005;
  reg n1009;
  wire [31:0] n1012;
  wire [31:0] n1014;
  wire n1016;
  wire n1029;
  wire n1031;
  wire n1035;
  wire [4:0] n1037;
  wire n1039;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1066;
  wire n1067;
  wire n1069;
  wire n1071;
  wire n1072;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1093;
  wire n1094;
  wire n1096;
  wire n1098;
  wire [15:0] n1099;
  reg n1103;
  wire [31:0] n1107;
  wire n1109;
  wire n1122;
  wire n1124;
  wire n1128;
  wire [4:0] n1130;
  wire n1132;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1159;
  wire n1160;
  wire n1162;
  wire n1164;
  wire n1165;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1186;
  wire n1187;
  wire n1189;
  wire n1191;
  wire [15:0] n1192;
  reg n1196;
  wire n1200;
  wire n1202;
  wire [3:0] n1205;
  wire [7:0] n1207;
  wire n1209;
  wire n1211;
  wire n1212;
  wire n1214;
  wire n1215;
  wire [7:0] n1216;
  wire n1218;
  wire n1220;
  wire [3:0] n1223;
  wire [3:0] n1224;
  wire n1226;
  wire [15:0] n1227;
  wire n1229;
  wire n1231;
  wire [3:0] n1234;
  wire [3:0] n1235;
  wire n1237;
  wire n1239;
  wire n1241;
  wire [3:0] n1244;
  wire [3:0] n1245;
  wire n1247;
  wire [2:0] n1249;
  reg [3:0] n1250;
  wire n1252;
  wire n1254;
  wire n1256;
  wire n1257;
  wire n1259;
  wire n1260;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1266;
  wire n1267;
  wire [30:0] n1268;
  wire [31:0] n1269;
  wire n1271;
  wire [30:0] n1272;
  wire [31:0] n1273;
  wire n1275;
  wire n1276;
  wire [2:0] n1279;
  wire [78:0] n1281;
  wire [79:0] n1283;
  wire n1285;
  wire n1287;
  wire [2:0] n1288;
  wire [79:0] n1289;
  wire n1292;
  wire [3:0] n1294;
  wire [7:0] n1296;
  wire n1298;
  wire [30:0] n1299;
  wire [31:0] n1300;
  wire n1302;
  wire [30:0] n1303;
  wire [31:0] n1304;
  wire n1306;
  wire n1307;
  wire [2:0] n1310;
  wire n1313;
  wire [2:0] n1316;
  wire [78:0] n1318;
  wire [79:0] n1319;
  wire n1321;
  wire n1323;
  wire [2:0] n1324;
  wire [79:0] n1325;
  wire n1328;
  wire [3:0] n1330;
  wire [7:0] n1332;
  wire n1334;
  wire [30:0] n1335;
  wire [31:0] n1336;
  wire n1338;
  wire [30:0] n1339;
  wire [31:0] n1340;
  wire n1342;
  wire n1343;
  wire [2:0] n1346;
  wire n1350;
  wire n1352;
  wire [2:0] n1353;
  wire [79:0] n1354;
  wire n1357;
  wire [3:0] n1359;
  wire [7:0] n1361;
  wire n1363;
  wire [6:0] n1365;
  wire n1367;
  wire [5:0] n1368;
  wire n1370;
  wire n1371;
  wire n1372;
  wire [5:0] n1373;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire [5:0] n1380;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire [5:0] n1386;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire [5:0] n1392;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire [5:0] n1398;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire [31:0] n1408;
  wire n1410;
  wire [4:0] n1411;
  reg [31:0] n1413;
  reg n1416;
  reg n1417;
  reg n1418;
  reg [2:0] n1419;
  reg [79:0] n1420;
  reg n1422;
  reg [3:0] n1425;
  reg [7:0] n1426;
  reg [6:0] n1427;
  reg n1429;
  wire n1431;
  wire n1433;
  wire n1434;
  wire [2:0] n1438;
  wire n1446;
  wire [14:0] n1448;
  wire [63:0] n1450;
  localparam [3:0] n1452 = 4'b0000;
  wire n1454;
  wire n1455;
  wire n1456;
  wire [62:0] n1457;
  wire n1459;
  wire n1460;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1470;
  wire n1472;
  wire n1473;
  wire [1:0] n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire [1:0] n1481;
  wire [1:0] n1482;
  wire [1:0] n1483;
  wire [1:0] n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1493;
  wire [3:0] n1494;
  wire [3:0] n1495;
  wire [3:0] n1496;
  wire [3:0] n1498;
  wire n1500;
  wire [7:0] n1501;
  wire n1503;
  wire [1:0] n1504;
  wire n1506;
  wire n1507;
  wire [4:0] n1508;
  wire n1510;
  wire n1511;
  wire [7:0] n1512;
  wire n1514;
  wire n1515;
  wire [7:0] n1516;
  wire n1517;
  wire n1519;
  wire n1521;
  wire n1523;
  wire n1525;
  wire n1532;
  wire n1534;
  wire n1536;
  wire n1538;
  wire n1540;
  wire n1543;
  wire [4:0] n1544;
  reg n1547;
  reg n1550;
  wire n1552;
  wire [5:0] n1553;
  reg n1559;
  reg n1565;
  wire n1567;
  wire [3:0] n1570;
  wire [7:0] n1572;
  wire n1574;
  wire [3:0] n1576;
  wire [7:0] n1577;
  wire n1578;
  wire [7:0] n1580;
  wire n1581;
  wire n1582;
  wire n1584;
  wire n1589;
  wire n1590;
  wire [31:0] n1592;
  wire [31:0] n1594;
  wire n1596;
  wire [3:0] n1599;
  wire [7:0] n1601;
  wire [5:0] n1603;
  wire [7:0] n1605;
  wire n1607;
  wire n1608;
  wire n1610;
  wire [3:0] n1613;
  wire [5:0] n1615;
  wire [7:0] n1617;
  wire [7:0] n1623;
  wire n1625;
  wire [2:0] n1626;
  wire n1628;
  wire [2:0] n1629;
  wire n1631;
  wire n1632;
  wire n1634;
  wire n1636;
  wire n1637;
  wire n1639;
  wire [3:0] n1642;
  wire n1644;
  wire [7:0] n1646;
  wire n1649;
  wire n1650;
  wire [3:0] n1652;
  wire n1653;
  wire n1654;
  wire n1656;
  wire n1657;
  wire [3:0] n1659;
  wire [7:0] n1661;
  wire n1663;
  wire [7:0] n1664;
  wire [2:0] n1665;
  wire n1667;
  wire [2:0] n1668;
  wire n1670;
  wire n1671;
  wire n1673;
  wire n1675;
  wire n1676;
  wire n1678;
  wire [3:0] n1681;
  wire n1683;
  wire [7:0] n1685;
  wire n1688;
  wire n1689;
  wire [3:0] n1691;
  wire n1692;
  wire n1693;
  wire n1695;
  wire n1696;
  wire [3:0] n1698;
  wire [7:0] n1700;
  wire n1702;
  wire [7:0] n1703;
  wire n1705;
  wire n1706;
  wire [3:0] n1708;
  wire n1709;
  wire n1710;
  wire [7:0] n1711;
  wire n1712;
  wire n1713;
  wire [3:0] n1714;
  wire [7:0] n1715;
  wire n1716;
  wire [7:0] n1717;
  wire n1719;
  wire [2:0] n1720;
  wire n1722;
  wire n1723;
  wire n1724;
  wire [2:0] n1725;
  wire n1727;
  wire n1729;
  wire n1731;
  wire [2:0] n1732;
  reg [31:0] n1734;
  wire [2:0] n1735;
  wire [1:0] n1743;
  wire n1745;
  wire [1:0] n1747;
  wire [1:0] n1748;
  wire [7:0] n1752;
  wire [31:0] n1754;
  wire n1756;
  wire n1765;
  wire n1767;
  wire [2:0] n1768;
  reg [31:0] n1769;
  reg [31:0] n1770;
  reg [31:0] n1771;
  wire [31:0] n1773;
  wire [31:0] n1774;
  wire [31:0] n1775;
  wire [31:0] n1776;
  wire [31:0] n1778;
  wire [31:0] n1779;
  wire [31:0] n1780;
  wire [31:0] n1781;
  wire n1783;
  wire n1785;
  wire n1787;
  wire n1788;
  wire n1790;
  wire n1791;
  wire n1793;
  wire n1794;
  wire n1796;
  wire n1797;
  wire n1799;
  wire n1800;
  wire n1802;
  wire n1803;
  wire n1805;
  wire n1806;
  wire n1808;
  wire n1809;
  wire n1811;
  wire n1812;
  wire n1814;
  wire n1815;
  wire n1817;
  wire n1818;
  wire n1820;
  wire n1821;
  wire n1823;
  wire n1824;
  wire n1826;
  wire n1827;
  wire n1829;
  wire n1830;
  wire n1832;
  wire n1833;
  wire n1835;
  wire n1836;
  wire n1838;
  wire n1839;
  wire n1841;
  wire n1842;
  wire n1844;
  wire n1845;
  wire n1847;
  wire n1848;
  wire n1850;
  wire n1851;
  wire n1853;
  wire n1854;
  wire n1856;
  wire n1857;
  wire n1859;
  wire n1860;
  wire n1862;
  wire n1863;
  wire n1865;
  wire n1866;
  wire n1868;
  wire n1869;
  wire n1871;
  wire n1872;
  wire n1874;
  wire n1875;
  wire n1877;
  wire n1878;
  wire n1880;
  wire n1881;
  wire n1883;
  wire n1884;
  wire n1886;
  wire n1887;
  wire n1889;
  wire n1890;
  wire n1892;
  wire n1893;
  wire n1895;
  wire n1896;
  wire n1898;
  wire n1899;
  wire n1927;
  wire [6:0] n1928;
  wire n1930;
  wire n1932;
  wire n1934;
  wire n1935;
  wire n1937;
  wire n1938;
  wire [3:0] n1941;
  wire [3:0] n1943;
  wire n1946;
  wire [3:0] n1948;
  wire n1950;
  wire [3:0] n1952;
  wire [6:0] n1953;
  wire n1955;
  wire n1957;
  wire n1959;
  wire [3:0] n1961;
  wire [7:0] n1963;
  wire n1964;
  wire n1965;
  wire n1967;
  wire [30:0] n1968;
  wire [31:0] n1969;
  wire n1971;
  wire n1973;
  wire [7:0] n1977;
  wire [2:0] n1980;
  wire [2:0] n1985;
  wire [6:0] n1987;
  wire [7:0] n1988;
  wire [8:0] n1990;
  wire [2:0] n1993;
  wire [22:0] n1995;
  wire [31:0] n1996;
  wire n1998;
  wire [2:0] n2001;
  wire [2:0] n2006;
  wire [10:0] n2009;
  wire [11:0] n2011;
  wire [2:0] n2014;
  wire [31:0] n2017;
  wire n2019;
  wire [2:0] n2037;
  wire [14:0] n2039;
  wire n2041;
  wire [2:0] n2044;
  wire [14:0] n2046;
  wire n2048;
  wire [2:0] n2051;
  wire [31:0] n2056;
  wire [2:0] n2059;
  wire [14:0] n2061;
  wire [30:0] n2062;
  wire [31:0] n2063;
  wire n2065;
  wire [2:0] n2068;
  wire [14:0] n2070;
  wire [30:0] n2071;
  wire [31:0] n2072;
  wire n2074;
  wire [2:0] n2077;
  wire [31:0] n2082;
  wire [2:0] n2085;
  wire [14:0] n2087;
  wire [30:0] n2088;
  wire [31:0] n2089;
  wire n2091;
  wire [2:0] n2094;
  wire [14:0] n2096;
  wire [30:0] n2097;
  wire [31:0] n2098;
  wire n2100;
  wire [2:0] n2103;
  wire [14:0] n2105;
  wire [30:0] n2106;
  wire [31:0] n2107;
  wire [31:0] n2109;
  wire [31:0] n2111;
  wire [5:0] n2112;
  wire [5:0] n2114;
  wire [5:0] n2116;
  wire [31:0] n2117;
  wire n2119;
  wire [2:0] n2122;
  wire [31:0] n2124;
  wire n2126;
  wire [2:0] n2129;
  wire [63:0] n2131;
  wire [30:0] n2132;
  wire [63:0] n2133;
  wire [31:0] n2134;
  wire n2137;
  wire n2138;
  wire n2139;
  wire [1:0] n2140;
  reg [31:0] n2142;
  wire [31:0] n2144;
  wire [2:0] n2147;
  wire [31:0] n2150;
  wire [31:0] n2152;
  wire [31:0] n2153;
  wire [31:0] n2154;
  wire [5:0] n2155;
  wire [31:0] n2156;
  wire [31:0] n2158;
  wire [5:0] n2159;
  wire [31:0] n2160;
  wire [31:0] n2161;
  wire [5:0] n2162;
  wire [31:0] n2163;
  wire [31:0] n2165;
  wire [5:0] n2166;
  wire [31:0] n2167;
  wire n2169;
  wire [2:0] n2172;
  wire n2177;
  wire [2:0] n2180;
  wire [3:0] n2184;
  reg [31:0] n2186;
  reg n2189;
  reg [2:0] n2192;
  reg [2:0] n2195;
  wire [79:0] n2196;
  reg [79:0] n2197;
  wire [15:0] n2198;
  reg [15:0] n2199;
  reg [5:0] n2203;
  reg [31:0] n2204;
  wire n2206;
  wire n2208;
  wire n2210;
  wire n2212;
  wire n2214;
  wire [3:0] n2215;
  reg n2217;
  reg [2:0] n2219;
  reg [2:0] n2221;
  wire n2223;
  wire [7:0] n2224;
  wire n2226;
  wire n2229;
  wire [3:0] n2232;
  wire n2234;
  wire n2236;
  wire [3:0] n2238;
  wire [7:0] n2240;
  wire n2242;
  wire n2243;
  wire [3:0] n2245;
  wire [7:0] n2246;
  wire n2247;
  wire [2:0] n2248;
  wire [2:0] n2249;
  wire [31:0] n2251;
  wire n2253;
  wire n2254;
  wire [3:0] n2256;
  wire [7:0] n2257;
  wire n2258;
  wire [2:0] n2259;
  wire [2:0] n2260;
  wire [95:0] n2261;
  wire [95:0] n2262;
  wire [5:0] n2266;
  wire [31:0] n2267;
  wire [31:0] n2269;
  wire n2270;
  wire n2271;
  wire [3:0] n2272;
  wire [7:0] n2273;
  wire n2274;
  wire [2:0] n2275;
  wire [2:0] n2276;
  wire [95:0] n2277;
  wire n2278;
  wire n2279;
  wire [5:0] n2283;
  wire [31:0] n2284;
  wire [31:0] n2285;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire [3:0] n2293;
  wire [7:0] n2294;
  wire n2295;
  wire [2:0] n2296;
  wire [2:0] n2297;
  wire [95:0] n2298;
  wire [6:0] n2299;
  wire n2300;
  wire [5:0] n2304;
  wire [31:0] n2305;
  wire [31:0] n2307;
  wire n2308;
  wire n2309;
  wire [31:0] n2310;
  wire [31:0] n2311;
  wire [31:0] n2312;
  wire [3:0] n2313;
  wire [7:0] n2314;
  wire n2315;
  wire [7:0] n2316;
  wire n2317;
  wire [2:0] n2318;
  wire [2:0] n2319;
  wire [95:0] n2320;
  wire [6:0] n2321;
  wire n2322;
  wire [5:0] n2326;
  wire [31:0] n2327;
  wire [31:0] n2329;
  wire n2331;
  wire n2332;
  wire [31:0] n2333;
  wire [31:0] n2334;
  wire [31:0] n2335;
  wire [3:0] n2336;
  wire [7:0] n2337;
  wire n2338;
  wire [5:0] n2339;
  wire [7:0] n2340;
  wire [7:0] n2343;
  wire n2344;
  wire [2:0] n2345;
  wire [2:0] n2346;
  wire [95:0] n2347;
  wire [6:0] n2348;
  wire n2349;
  wire [5:0] n2353;
  wire [31:0] n2354;
  wire [31:0] n2355;
  wire n2357;
  wire n2358;
  wire [31:0] n2359;
  wire [31:0] n2360;
  wire [31:0] n2361;
  wire [3:0] n2362;
  wire [7:0] n2364;
  wire [7:0] n2365;
  wire n2366;
  wire [5:0] n2367;
  wire [7:0] n2368;
  wire [7:0] n2371;
  wire n2372;
  wire [2:0] n2373;
  wire [2:0] n2374;
  wire [95:0] n2375;
  wire [6:0] n2376;
  wire n2377;
  wire [5:0] n2381;
  wire [31:0] n2382;
  wire [31:0] n2384;
  wire n2386;
  wire n2387;
  wire [31:0] n2388;
  wire [31:0] n2389;
  wire [31:0] n2390;
  wire [3:0] n2392;
  wire [7:0] n2394;
  wire [7:0] n2395;
  wire n2396;
  wire [5:0] n2397;
  wire [7:0] n2398;
  wire [7:0] n2401;
  wire n2402;
  wire [2:0] n2403;
  wire [2:0] n2404;
  wire [95:0] n2405;
  wire [6:0] n2406;
  wire n2407;
  wire [5:0] n2411;
  wire [31:0] n2412;
  wire [31:0] n2414;
  wire n2416;
  wire n2417;
  wire [31:0] n2418;
  wire [31:0] n2419;
  wire [31:0] n2420;
  wire [3:0] n2421;
  wire [7:0] n2423;
  wire [7:0] n2424;
  wire n2425;
  wire [5:0] n2426;
  wire [7:0] n2427;
  wire [7:0] n2430;
  wire n2431;
  wire [2:0] n2432;
  wire [2:0] n2433;
  wire [95:0] n2434;
  wire [6:0] n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire [5:0] n2442;
  wire [31:0] n2443;
  wire [31:0] n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire [2:0] n2448;
  wire [79:0] n2449;
  wire n2451;
  wire [31:0] n2452;
  wire [27:0] n2453;
  wire [27:0] n2454;
  wire [27:0] n2455;
  wire [3:0] n2456;
  wire [3:0] n2457;
  wire [31:0] n2458;
  wire [3:0] n2459;
  wire [7:0] n2461;
  wire [7:0] n2462;
  wire n2463;
  wire [5:0] n2464;
  wire [7:0] n2465;
  wire [7:0] n2468;
  wire n2469;
  wire [2:0] n2470;
  wire [2:0] n2471;
  wire [95:0] n2472;
  wire [6:0] n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire [5:0] n2480;
  wire [31:0] n2481;
  wire [31:0] n2483;
  wire n2485;
  wire n2486;
  wire n2487;
  wire [2:0] n2488;
  wire [79:0] n2489;
  wire n2491;
  wire [31:0] n2492;
  wire [31:0] n2493;
  wire [27:0] n2494;
  wire [27:0] n2495;
  wire [27:0] n2496;
  wire [3:0] n2497;
  wire [3:0] n2498;
  wire [31:0] n2499;
  wire [3:0] n2501;
  wire [7:0] n2503;
  wire [7:0] n2504;
  wire n2505;
  wire [5:0] n2506;
  wire [7:0] n2507;
  wire [7:0] n2510;
  wire n2511;
  wire [2:0] n2512;
  wire [2:0] n2513;
  wire [95:0] n2514;
  wire [6:0] n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire [5:0] n2522;
  wire [31:0] n2523;
  wire [31:0] n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire [2:0] n2529;
  wire [79:0] n2530;
  wire n2532;
  wire [31:0] n2533;
  wire [31:0] n2534;
  wire [31:0] n2535;
  wire [31:0] n2536;
  wire [3:0] n2537;
  wire [7:0] n2539;
  wire [7:0] n2540;
  wire n2541;
  wire [5:0] n2542;
  wire [7:0] n2543;
  wire [7:0] n2546;
  wire n2547;
  wire [2:0] n2548;
  wire [2:0] n2549;
  wire [95:0] n2550;
  wire [6:0] n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire [5:0] n2558;
  wire [31:0] n2559;
  wire [31:0] n2560;
  wire n2562;
  wire n2563;
  wire n2564;
  wire [2:0] n2565;
  wire [79:0] n2566;
  wire n2568;
  wire [31:0] n2569;
  wire [31:0] n2570;
  wire [31:0] n2571;
  wire [3:0] n2573;
  wire [7:0] n2575;
  wire [7:0] n2576;
  wire n2577;
  wire [5:0] n2578;
  wire [7:0] n2579;
  wire [7:0] n2582;
  wire n2583;
  wire [2:0] n2584;
  wire [2:0] n2585;
  wire [95:0] n2586;
  wire [6:0] n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire [5:0] n2594;
  wire [31:0] n2595;
  wire [31:0] n2596;
  wire n2598;
  wire n2599;
  wire n2600;
  wire [2:0] n2601;
  wire [79:0] n2602;
  wire n2604;
  wire [31:0] n2605;
  wire [31:0] n2606;
  wire [31:0] n2607;
  wire [3:0] n2609;
  wire [7:0] n2611;
  wire [7:0] n2612;
  wire n2613;
  wire [5:0] n2614;
  wire [7:0] n2615;
  wire [7:0] n2618;
  wire n2619;
  wire [2:0] n2620;
  wire [2:0] n2621;
  wire [95:0] n2622;
  wire [6:0] n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire [5:0] n2630;
  wire [31:0] n2631;
  wire [31:0] n2633;
  wire n2635;
  wire n2637;
  wire n2638;
  wire [2:0] n2639;
  wire [79:0] n2640;
  wire n2642;
  wire [31:0] n2643;
  wire [31:0] n2644;
  wire [31:0] n2645;
  wire [3:0] n2647;
  wire [7:0] n2649;
  wire [7:0] n2650;
  wire n2651;
  wire [5:0] n2652;
  wire [7:0] n2653;
  wire [7:0] n2657;
  wire n2658;
  wire [2:0] n2659;
  wire [2:0] n2660;
  wire [95:0] n2661;
  wire [6:0] n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire [5:0] n2669;
  wire [31:0] n2670;
  wire [31:0] n2672;
  wire n2674;
  wire n2676;
  wire n2677;
  wire [2:0] n2678;
  wire [79:0] n2679;
  wire n2681;
  wire [31:0] n2682;
  wire [31:0] n2683;
  wire [31:0] n2684;
  wire [3:0] n2686;
  wire [7:0] n2688;
  wire [7:0] n2689;
  wire n2690;
  wire [5:0] n2691;
  wire [7:0] n2692;
  wire [7:0] n2696;
  wire n2697;
  wire [2:0] n2698;
  wire [2:0] n2699;
  wire [95:0] n2700;
  wire [6:0] n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire [5:0] n2708;
  wire [31:0] n2709;
  wire [31:0] n2711;
  wire n2713;
  wire n2715;
  wire n2716;
  wire [2:0] n2717;
  wire [79:0] n2718;
  wire n2720;
  wire [31:0] n2721;
  wire [31:0] n2722;
  wire [31:0] n2723;
  wire [3:0] n2725;
  wire [7:0] n2727;
  wire [7:0] n2728;
  wire n2729;
  wire [5:0] n2730;
  wire [7:0] n2731;
  wire [7:0] n2735;
  wire n2736;
  wire [2:0] n2737;
  wire [2:0] n2738;
  wire [95:0] n2739;
  wire [6:0] n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire [5:0] n2747;
  wire [31:0] n2748;
  wire [31:0] n2750;
  wire n2753;
  wire n2755;
  wire n2756;
  wire [2:0] n2757;
  wire [79:0] n2758;
  wire n2760;
  wire [31:0] n2761;
  wire [31:0] n2762;
  wire [31:0] n2763;
  wire [15:0] n2764;
  wire [31:0] n2765;
  wire [3:0] n2766;
  wire [7:0] n2768;
  wire [7:0] n2769;
  wire n2770;
  wire [5:0] n2771;
  wire [7:0] n2772;
  wire [7:0] n2775;
  wire n2776;
  wire [2:0] n2777;
  wire [2:0] n2778;
  wire [95:0] n2779;
  wire [6:0] n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire [5:0] n2787;
  wire [31:0] n2788;
  wire n2790;
  wire n2792;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2798;
  wire n2799;
  wire [7:0] n2800;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire [6:0] n2806;
  wire [23:0] n2808;
  wire [79:0] n2810;
  wire n2811;
  wire [5:0] n2812;
  wire [22:0] n2814;
  wire [23:0] n2816;
  wire [79:0] n2818;
  wire n2819;
  wire [4:0] n2820;
  wire [21:0] n2822;
  wire [23:0] n2824;
  wire [79:0] n2826;
  wire n2827;
  wire [3:0] n2828;
  wire [20:0] n2830;
  wire [23:0] n2832;
  wire [79:0] n2834;
  wire n2835;
  wire [2:0] n2836;
  wire [19:0] n2838;
  wire [23:0] n2840;
  wire [79:0] n2842;
  wire n2843;
  wire [1:0] n2844;
  wire [18:0] n2846;
  wire [23:0] n2848;
  wire [79:0] n2850;
  wire n2851;
  wire [17:0] n2853;
  wire [23:0] n2855;
  wire [79:0] n2857;
  wire [79:0] n2858;
  wire [79:0] n2859;
  wire [79:0] n2860;
  wire [79:0] n2861;
  wire [79:0] n2862;
  wire [79:0] n2863;
  wire [7:0] n2864;
  wire n2866;
  wire [7:0] n2867;
  wire [7:0] n2868;
  wire [7:0] n2870;
  wire [24:0] n2872;
  wire [79:0] n2874;
  wire [79:0] n2876;
  wire [79:0] n2877;
  wire [79:0] n2879;
  wire n2881;
  wire n2883;
  wire n2884;
  wire n2885;
  wire [31:0] n2887;
  wire [79:0] n2889;
  wire [15:0] n2890;
  wire [15:0] n2892;
  wire [31:0] n2894;
  wire [79:0] n2896;
  wire [79:0] n2897;
  wire [79:0] n2899;
  wire n2901;
  wire [32:0] n2903;
  wire [79:0] n2905;
  wire n2907;
  wire [2:0] n2908;
  reg [79:0] n2910;
  wire n2912;
  wire n2914;
  wire n2915;
  wire [30:0] n2916;
  wire [31:0] n2917;
  wire n2919;
  wire [2:0] n2922;
  wire n2926;
  wire [3:0] n2928;
  wire [7:0] n2930;
  wire [79:0] n2931;
  wire n2933;
  wire [7:0] n2934;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire [6:0] n2940;
  wire [23:0] n2942;
  wire [79:0] n2944;
  wire n2945;
  wire [5:0] n2946;
  wire [22:0] n2948;
  wire [23:0] n2950;
  wire [79:0] n2952;
  wire n2953;
  wire [4:0] n2954;
  wire [21:0] n2956;
  wire [23:0] n2958;
  wire [79:0] n2960;
  wire n2961;
  wire [3:0] n2962;
  wire [20:0] n2964;
  wire [23:0] n2966;
  wire [79:0] n2968;
  wire n2969;
  wire [2:0] n2970;
  wire [19:0] n2972;
  wire [23:0] n2974;
  wire [79:0] n2976;
  wire n2977;
  wire [1:0] n2978;
  wire [18:0] n2980;
  wire [23:0] n2982;
  wire [79:0] n2984;
  wire n2985;
  wire [17:0] n2987;
  wire [23:0] n2989;
  wire [79:0] n2991;
  wire [79:0] n2992;
  wire [79:0] n2993;
  wire [79:0] n2994;
  wire [79:0] n2995;
  wire [79:0] n2996;
  wire [79:0] n2997;
  wire [7:0] n2998;
  wire n3000;
  wire [7:0] n3001;
  wire [7:0] n3002;
  wire [7:0] n3004;
  wire [24:0] n3006;
  wire [79:0] n3008;
  wire [79:0] n3010;
  wire [79:0] n3011;
  wire [79:0] n3013;
  wire n3015;
  wire [15:0] n3016;
  wire n3018;
  wire n3019;
  wire n3020;
  wire [15:0] n3021;
  wire [31:0] n3023;
  wire [79:0] n3025;
  wire [15:0] n3026;
  wire [15:0] n3027;
  wire [15:0] n3029;
  wire [31:0] n3031;
  wire [79:0] n3033;
  wire [79:0] n3034;
  wire [79:0] n3036;
  wire n3038;
  wire n3040;
  wire n3041;
  wire n3042;
  wire [47:0] n3044;
  wire [79:0] n3046;
  wire [31:0] n3047;
  wire [31:0] n3049;
  wire [47:0] n3051;
  wire [79:0] n3053;
  wire [79:0] n3054;
  wire [79:0] n3056;
  wire n3058;
  wire [2:0] n3059;
  reg [79:0] n3061;
  wire n3063;
  wire n3065;
  wire n3067;
  wire n3069;
  wire n3071;
  wire n3073;
  wire n3075;
  wire n3077;
  wire n3079;
  wire n3081;
  wire n3083;
  wire [7:0] n3084;
  wire n3086;
  wire n3087;
  wire n3088;
  wire [7:0] n3089;
  wire [24:0] n3091;
  wire [76:0] n3093;
  wire [79:0] n3095;
  wire [7:0] n3096;
  wire [7:0] n3097;
  wire [24:0] n3099;
  wire [24:0] n3101;
  wire [76:0] n3103;
  wire [79:0] n3105;
  wire [79:0] n3106;
  wire [79:0] n3108;
  wire n3110;
  wire [15:0] n3111;
  wire n3113;
  wire n3114;
  wire n3115;
  wire [15:0] n3116;
  wire [32:0] n3118;
  wire [76:0] n3120;
  wire [79:0] n3122;
  wire [15:0] n3123;
  wire [15:0] n3124;
  wire [32:0] n3126;
  wire [32:0] n3128;
  wire [76:0] n3130;
  wire [79:0] n3132;
  wire [79:0] n3133;
  wire [79:0] n3135;
  wire n3137;
  wire n3139;
  wire n3140;
  wire n3141;
  wire [48:0] n3143;
  wire [76:0] n3145;
  wire [79:0] n3147;
  wire [31:0] n3148;
  wire [48:0] n3150;
  wire [48:0] n3152;
  wire [76:0] n3154;
  wire [79:0] n3156;
  wire [79:0] n3157;
  wire [79:0] n3159;
  wire n3161;
  wire [7:0] n3162;
  wire n3164;
  wire [22:0] n3165;
  wire n3167;
  wire n3168;
  wire [15:0] n3170;
  wire [79:0] n3172;
  wire n3173;
  wire [16:0] n3175;
  wire [17:0] n3177;
  wire [22:0] n3178;
  wire [40:0] n3179;
  wire [76:0] n3181;
  wire [79:0] n3183;
  wire [79:0] n3184;
  wire [7:0] n3185;
  wire n3187;
  wire [22:0] n3188;
  wire n3190;
  wire n3191;
  wire [15:0] n3193;
  wire [79:0] n3195;
  wire n3196;
  wire [15:0] n3198;
  wire [16:0] n3200;
  wire [22:0] n3201;
  wire [39:0] n3202;
  wire [79:0] n3204;
  wire [79:0] n3205;
  wire n3206;
  wire [15:0] n3208;
  wire [16:0] n3210;
  wire [22:0] n3211;
  wire [39:0] n3212;
  wire [79:0] n3214;
  wire [79:0] n3215;
  wire [79:0] n3216;
  wire n3218;
  wire [10:0] n3219;
  wire n3221;
  wire n3222;
  wire [15:0] n3224;
  wire [79:0] n3226;
  wire [10:0] n3227;
  wire n3229;
  wire n3230;
  wire [15:0] n3232;
  wire [19:0] n3233;
  wire [35:0] n3234;
  wire [79:0] n3236;
  wire n3237;
  wire [15:0] n3239;
  wire [16:0] n3241;
  wire [19:0] n3242;
  wire [36:0] n3243;
  wire [79:0] n3245;
  wire [79:0] n3246;
  wire [79:0] n3247;
  wire n3249;
  wire [4:0] n3250;
  reg [79:0] n3252;
  wire n3255;
  wire n3257;
  wire n3259;
  wire n3261;
  wire [7:0] n3262;
  reg [3:0] n3272;
  reg n3276;
  reg [6:0] n3277;
  reg [79:0] n3279;
  wire n3281;
  wire [7:0] n3282;
  reg [3:0] n3289;
  reg n3292;
  reg [6:0] n3293;
  reg [79:0] n3297;
  wire [3:0] n3298;
  wire n3300;
  wire [6:0] n3301;
  wire [79:0] n3302;
  wire n3304;
  wire n3306;
  wire n3307;
  wire n3309;
  wire n3310;
  wire n3317;
  wire [14:0] n3319;
  wire [63:0] n3321;
  localparam [3:0] n3323 = 4'b0000;
  wire n3325;
  wire n3326;
  wire n3327;
  wire [62:0] n3328;
  wire n3330;
  wire n3331;
  wire n3334;
  wire n3335;
  wire n3336;
  wire n3337;
  wire n3338;
  wire n3339;
  wire n3341;
  wire n3343;
  wire n3344;
  wire [1:0] n3346;
  wire n3347;
  wire n3348;
  wire n3349;
  wire n3350;
  wire n3351;
  wire [1:0] n3352;
  wire [1:0] n3353;
  wire [1:0] n3354;
  wire [1:0] n3355;
  wire n3356;
  wire n3357;
  wire n3358;
  wire n3359;
  wire n3360;
  wire n3364;
  wire n3366;
  wire n3373;
  wire [14:0] n3375;
  wire [63:0] n3377;
  localparam [3:0] n3379 = 4'b0000;
  wire n3381;
  wire n3382;
  wire n3383;
  wire [62:0] n3384;
  wire n3386;
  wire n3387;
  wire n3390;
  wire n3391;
  wire n3392;
  wire n3393;
  wire n3394;
  wire n3395;
  wire n3397;
  wire n3399;
  wire n3400;
  wire [1:0] n3402;
  wire n3403;
  wire n3404;
  wire n3405;
  wire n3406;
  wire n3407;
  wire [1:0] n3408;
  wire [1:0] n3409;
  wire [1:0] n3410;
  wire [1:0] n3411;
  wire n3412;
  wire n3413;
  wire n3414;
  wire n3415;
  wire n3416;
  wire n3420;
  wire n3422;
  wire n3423;
  wire n3425;
  wire n3426;
  wire n3428;
  wire n3429;
  wire n3431;
  wire n3432;
  wire n3434;
  wire n3435;
  wire n3437;
  wire n3438;
  wire n3440;
  wire n3441;
  wire n3443;
  wire n3444;
  wire n3446;
  wire n3447;
  wire n3449;
  wire n3450;
  wire n3452;
  wire n3453;
  wire n3455;
  wire n3456;
  wire n3458;
  wire n3459;
  wire n3461;
  wire n3462;
  wire n3464;
  wire n3465;
  wire n3467;
  wire n3468;
  wire n3470;
  wire n3471;
  wire n3473;
  wire n3474;
  wire [14:0] n3475;
  wire n3477;
  wire n3478;
  wire [62:0] n3479;
  wire n3481;
  wire n3482;
  wire n3483;
  wire [62:0] n3484;
  wire n3486;
  wire n3487;
  wire n3489;
  wire n3491;
  wire n3492;
  wire n3494;
  wire n3495;
  wire n3496;
  wire n3497;
  wire [79:0] n3499;
  wire n3501;
  wire n3503;
  wire n3504;
  wire n3506;
  wire n3507;
  wire [1:0] n3508;
  reg [3:0] n3510;
  reg n3512;
  reg [6:0] n3513;
  reg [79:0] n3514;
  reg [79:0] n3516;
  wire [3:0] n3518;
  wire n3520;
  wire [6:0] n3521;
  wire [79:0] n3522;
  wire [79:0] n3523;
  wire [3:0] n3525;
  wire n3526;
  wire [6:0] n3527;
  wire [79:0] n3528;
  wire [79:0] n3529;
  wire n3530;
  wire n3531;
  wire n3533;
  wire [3:0] n3536;
  wire [7:0] n3538;
  wire n3540;
  wire n3541;
  wire [3:0] n3543;
  wire [7:0] n3544;
  wire n3546;
  wire n3547;
  wire [3:0] n3548;
  wire [7:0] n3549;
  wire n3550;
  wire [6:0] n3551;
  wire [79:0] n3552;
  wire [79:0] n3553;
  wire n3554;
  wire n3555;
  wire n3557;
  wire [7:0] n3561;
  wire n3562;
  wire [7:0] n3564;
  wire n3565;
  wire [3:0] n3567;
  wire [7:0] n3568;
  wire n3570;
  wire [6:0] n3571;
  wire n3572;
  wire [6:0] n3573;
  wire [79:0] n3574;
  wire n3575;
  wire n3576;
  wire [3:0] n3577;
  wire [3:0] n3578;
  wire [3:0] n3579;
  wire [3:0] n3581;
  wire [7:0] n3582;
  wire n3583;
  wire [6:0] n3584;
  wire n3585;
  wire [6:0] n3586;
  wire [79:0] n3587;
  wire [79:0] n3588;
  wire n3589;
  wire n3591;
  wire [3:0] n3592;
  wire [7:0] n3593;
  wire n3594;
  wire [6:0] n3595;
  wire n3596;
  wire [6:0] n3597;
  wire [79:0] n3598;
  wire [79:0] n3599;
  wire n3600;
  wire [3:0] n3601;
  wire [3:0] n3602;
  wire [3:0] n3604;
  wire [7:0] n3605;
  wire n3606;
  wire [6:0] n3607;
  wire n3608;
  wire [6:0] n3609;
  wire [79:0] n3610;
  wire [79:0] n3611;
  wire n3612;
  wire [3:0] n3613;
  wire [3:0] n3614;
  wire [3:0] n3615;
  wire [7:0] n3616;
  wire n3618;
  wire [6:0] n3619;
  wire [79:0] n3620;
  wire [79:0] n3621;
  wire n3622;
  wire [6:0] n3623;
  wire [79:0] n3624;
  wire [79:0] n3625;
  wire n3626;
  wire [3:0] n3627;
  wire [3:0] n3628;
  wire [3:0] n3630;
  wire [7:0] n3631;
  wire n3633;
  wire [6:0] n3635;
  wire [79:0] n3636;
  wire [79:0] n3637;
  wire n3638;
  wire [6:0] n3639;
  wire [79:0] n3640;
  wire [79:0] n3641;
  wire n3643;
  wire [31:0] n3644;
  wire n3646;
  wire [31:0] n3647;
  wire [31:0] n3649;
  wire [7:0] n3650;
  wire [7:0] n3651;
  wire n3652;
  wire n3654;
  wire n3656;
  wire [3:0] n3658;
  wire [7:0] n3660;
  wire n3661;
  wire [1:0] n3662;
  wire [1:0] n3663;
  wire n3667;
  wire n3668;
  wire n3669;
  wire n3670;
  wire n3672;
  wire n3674;
  wire [3:0] n3676;
  wire [7:0] n3678;
  wire n3679;
  wire [1:0] n3680;
  wire [1:0] n3681;
  wire n3685;
  wire n3686;
  wire n3687;
  wire n3689;
  wire n3691;
  wire n3692;
  wire n3694;
  wire [31:0] n3695;
  wire n3697;
  wire n3699;
  wire [3:0] n3701;
  wire n3702;
  wire n3703;
  wire n3704;
  wire n3705;
  wire [79:0] n3706;
  wire n3707;
  wire n3708;
  wire n3709;
  wire n3710;
  wire n3712;
  wire n3714;
  wire n3715;
  wire [7:0] n3716;
  wire [7:0] n3717;
  wire [7:0] n3718;
  wire [15:0] n3719;
  wire [1:0] n3730;
  wire n3732;
  wire n3736;
  wire n3742;
  wire [15:0] n3743;
  wire n3745;
  wire [5:0] n3746;
  wire n3748;
  wire n3749;
  wire n3752;
  wire n3755;
  wire n3756;
  wire n3758;
  wire n3759;
  wire n3761;
  wire n3767;
  wire [1:0] n3768;
  wire n3770;
  wire n3771;
  wire [1:0] n3772;
  wire [1:0] n3774;
  wire n3776;
  wire [14:0] n3777;
  wire n3779;
  wire [14:0] n3780;
  wire n3782;
  wire n3783;
  wire [15:0] n3785;
  wire [16:0] n3787;
  wire [22:0] n3788;
  wire [39:0] n3789;
  wire [79:0] n3791;
  wire [79:0] n3792;
  wire [79:0] n3794;
  wire n3796;
  wire [14:0] n3797;
  wire n3799;
  wire [14:0] n3800;
  wire n3802;
  wire n3803;
  wire [15:0] n3805;
  wire [63:0] n3806;
  wire [79:0] n3807;
  wire [79:0] n3808;
  wire [79:0] n3810;
  wire n3812;
  wire [2:0] n3813;
  reg n3815;
  reg [79:0] n3816;
  wire n3817;
  wire [1:0] n3818;
  wire [79:0] n3819;
  wire n3821;
  wire n3822;
  wire [1:0] n3823;
  wire [3:0] n3826;
  wire [7:0] n3827;
  wire [79:0] n3828;
  wire [31:0] n3829;
  wire n3831;
  wire n3833;
  wire n3835;
  wire n3836;
  wire n3838;
  wire n3839;
  wire n3841;
  wire n3843;
  wire [78:0] n3844;
  wire [79:0] n3846;
  wire n3848;
  wire n3849;
  wire n3850;
  wire [78:0] n3851;
  wire [79:0] n3852;
  wire [79:0] n3853;
  wire [79:0] n3854;
  wire [79:0] n3855;
  wire n3857;
  wire n3859;
  wire n3866;
  wire [14:0] n3868;
  wire [63:0] n3870;
  localparam [3:0] n3872 = 4'b0000;
  wire n3874;
  wire n3875;
  wire n3876;
  wire [62:0] n3877;
  wire n3879;
  wire n3880;
  wire n3883;
  wire n3884;
  wire n3885;
  wire n3886;
  wire n3887;
  wire n3888;
  wire n3890;
  wire n3892;
  wire n3893;
  wire [1:0] n3895;
  wire n3896;
  wire n3897;
  wire n3898;
  wire n3899;
  wire n3900;
  wire [1:0] n3901;
  wire [1:0] n3902;
  wire [1:0] n3903;
  wire [1:0] n3904;
  wire n3905;
  wire n3906;
  wire n3907;
  wire n3908;
  wire n3909;
  wire n3918;
  wire [14:0] n3920;
  wire [63:0] n3922;
  localparam [3:0] n3924 = 4'b0000;
  wire n3926;
  wire n3927;
  wire n3928;
  wire [62:0] n3929;
  wire n3931;
  wire n3932;
  wire n3935;
  wire n3936;
  wire n3937;
  wire n3938;
  wire n3939;
  wire n3940;
  wire n3942;
  wire n3944;
  wire n3945;
  wire [1:0] n3947;
  wire n3948;
  wire n3949;
  wire n3950;
  wire n3951;
  wire n3952;
  wire [1:0] n3953;
  wire [1:0] n3954;
  wire [1:0] n3955;
  wire [1:0] n3956;
  wire n3957;
  wire n3958;
  wire n3959;
  wire n3960;
  wire n3961;
  wire [3:0] n3964;
  wire [3:0] n3965;
  wire [3:0] n3966;
  wire n3968;
  wire [3:0] n3969;
  wire [3:0] n3970;
  wire [3:0] n3973;
  wire [7:0] n3975;
  wire n3976;
  wire [3:0] n3977;
  wire [3:0] n3978;
  wire [3:0] n3980;
  wire [7:0] n3981;
  wire [79:0] n3982;
  wire n3983;
  wire [3:0] n3984;
  wire [3:0] n3985;
  wire [3:0] n3986;
  wire [7:0] n3988;
  wire [7:0] n3989;
  wire n3990;
  wire n3991;
  wire [31:0] n3992;
  wire [27:0] n3993;
  wire [27:0] n3994;
  wire [27:0] n3995;
  wire [3:0] n3996;
  wire [3:0] n3997;
  wire n3998;
  wire [1:0] n3999;
  wire [3:0] n4000;
  wire [7:0] n4002;
  wire [7:0] n4003;
  wire [79:0] n4004;
  wire n4005;
  wire n4006;
  wire n4007;
  wire n4008;
  wire [79:0] n4009;
  wire n4010;
  wire n4011;
  wire [31:0] n4012;
  wire [31:0] n4013;
  wire n4014;
  wire [1:0] n4015;
  wire [3:0] n4016;
  wire [7:0] n4017;
  wire [7:0] n4018;
  wire [79:0] n4019;
  wire n4020;
  wire n4021;
  wire n4022;
  wire n4023;
  wire [79:0] n4024;
  wire n4026;
  wire n4027;
  wire [31:0] n4028;
  wire n4029;
  wire [1:0] n4030;
  wire [3:0] n4032;
  wire [7:0] n4034;
  wire [7:0] n4035;
  wire [79:0] n4036;
  wire n4037;
  wire n4038;
  wire n4039;
  wire n4040;
  wire [79:0] n4041;
  wire n4043;
  wire n4045;
  wire n4047;
  wire n4049;
  wire [30:0] n4050;
  wire [31:0] n4051;
  wire n4053;
  wire n4055;
  wire n4057;
  wire [2:0] n4058;
  wire [79:0] n4059;
  wire n4061;
  wire [7:0] n4065;
  wire n4067;
  wire n4068;
  wire n4069;
  wire n4070;
  wire n4071;
  wire n4072;
  wire [3:0] n4074;
  wire [7:0] n4075;
  wire n4077;
  wire n4079;
  wire [30:0] n4080;
  wire [31:0] n4081;
  wire n4083;
  wire n4091;
  wire [2:0] n4092;
  wire [79:0] n4093;
  wire n4095;
  wire [2:0] n4096;
  wire [30:0] n4097;
  wire [31:0] n4098;
  wire n4100;
  wire [14:0] n4101;
  wire n4103;
  wire [2:0] n4104;
  wire [14:0] n4111;
  wire n4113;
  wire [2:0] n4114;
  wire [14:0] n4121;
  wire n4123;
  wire [2:0] n4124;
  wire [14:0] n4131;
  wire n4133;
  wire [2:0] n4134;
  wire [14:0] n4141;
  wire n4143;
  wire [2:0] n4144;
  wire [2:0] n4151;
  wire [2:0] n4160;
  wire [79:0] n4163;
  wire [2:0] n4166;
  wire [79:0] n4168;
  wire [2:0] n4171;
  wire [79:0] n4173;
  wire [2:0] n4176;
  wire [79:0] n4178;
  wire [2:0] n4181;
  wire [79:0] n4182;
  wire n4186;
  wire [2:0] n4187;
  wire [79:0] n4188;
  wire n4190;
  wire n4192;
  wire n4194;
  wire n4195;
  wire [30:0] n4196;
  wire [31:0] n4197;
  wire n4199;
  wire n4207;
  wire [2:0] n4208;
  wire [79:0] n4209;
  wire n4211;
  wire n4214;
  wire n4215;
  wire n4216;
  wire n4217;
  wire n4220;
  wire [2:0] n4221;
  wire [79:0] n4222;
  wire n4223;
  wire n4230;
  wire [14:0] n4232;
  wire [63:0] n4234;
  localparam [3:0] n4236 = 4'b0000;
  wire n4238;
  wire n4239;
  wire n4240;
  wire [62:0] n4241;
  wire n4243;
  wire n4244;
  wire n4247;
  wire n4248;
  wire n4249;
  wire n4250;
  wire n4251;
  wire n4252;
  wire n4254;
  wire n4256;
  wire n4257;
  wire [1:0] n4259;
  wire n4260;
  wire n4261;
  wire n4262;
  wire n4263;
  wire n4264;
  wire [1:0] n4265;
  wire [1:0] n4266;
  wire [1:0] n4267;
  wire [1:0] n4268;
  wire n4269;
  wire n4270;
  wire n4271;
  wire n4272;
  wire n4273;
  wire n4278;
  wire n4279;
  wire n4280;
  wire n4281;
  wire n4284;
  wire n4285;
  wire n4286;
  wire n4287;
  wire n4290;
  wire n4291;
  wire n4292;
  wire n4293;
  wire n4296;
  wire n4297;
  wire n4298;
  wire n4299;
  wire n4302;
  wire n4303;
  wire n4304;
  wire n4305;
  wire n4307;
  wire n4309;
  wire n4310;
  wire [6:0] n4311;
  wire [2:0] n4312;
  wire [6:0] n4313;
  wire [6:0] n4314;
  wire n4316;
  wire n4318;
  wire n4319;
  wire [31:0] n4320;
  wire n4322;
  wire [31:0] n4323;
  wire [31:0] n4325;
  wire [31:0] n4326;
  wire [31:0] n4327;
  wire n4329;
  wire n4330;
  wire n4333;
  wire [2:0] n4334;
  wire [79:0] n4335;
  wire n4336;
  wire [12:0] n4337;
  wire [3:0] n4338;
  wire [12:0] n4339;
  wire [12:0] n4340;
  wire [3:0] n4341;
  wire [3:0] n4342;
  wire [3:0] n4344;
  wire n4345;
  wire n4346;
  wire n4348;
  wire n4350;
  wire n4353;
  wire n4357;
  wire n4361;
  wire n4365;
  wire n4369;
  wire n4373;
  wire n4377;
  wire n4381;
  wire [7:0] n4383;
  wire n4384;
  reg n4385;
  wire n4386;
  reg n4387;
  wire n4388;
  reg n4389;
  wire n4390;
  reg n4391;
  wire n4392;
  reg n4393;
  wire n4394;
  reg n4395;
  wire n4396;
  reg n4397;
  wire n4398;
  reg n4399;
  wire n4400;
  reg n4401;
  wire n4402;
  reg n4403;
  wire n4404;
  reg n4405;
  wire n4406;
  reg n4407;
  wire n4408;
  wire n4411;
  wire n4413;
  wire n4414;
  wire n4417;
  wire n4419;
  wire n4420;
  wire n4423;
  wire n4425;
  wire n4426;
  wire n4429;
  wire n4431;
  wire n4432;
  wire n4435;
  wire n4437;
  wire n4438;
  wire n4441;
  wire n4443;
  wire [5:0] n4444;
  reg n4446;
  wire n4448;
  wire [31:0] n4450;
  wire n4452;
  wire n4454;
  wire [31:0] n4456;
  wire n4458;
  wire n4460;
  wire n4462;
  wire n4463;
  wire [31:0] n4465;
  wire n4467;
  wire n4469;
  wire n4471;
  wire n4472;
  wire [31:0] n4474;
  wire n4476;
  wire n4479;
  wire n4480;
  wire n4481;
  wire n4483;
  wire [31:0] n4484;
  wire [31:0] n4486;
  wire [2:0] n4487;
  wire [2:0] n4489;
  wire [31:0] n4491;
  wire [31:0] n4493;
  wire n4496;
  wire n4497;
  wire n4498;
  wire n4500;
  wire [31:0] n4501;
  wire [31:0] n4503;
  wire [2:0] n4504;
  wire [2:0] n4506;
  wire [31:0] n4508;
  wire [31:0] n4510;
  wire n4513;
  wire n4514;
  wire n4515;
  wire n4517;
  wire [31:0] n4518;
  wire [31:0] n4520;
  wire [2:0] n4521;
  wire [2:0] n4523;
  wire [31:0] n4527;
  wire [31:0] n4529;
  wire n4532;
  wire n4533;
  wire n4534;
  wire n4539;
  wire n4540;
  wire n4541;
  wire [8:0] n4542;
  reg [31:0] n4546;
  wire [31:0] n4547;
  wire [31:0] n4548;
  wire n4550;
  wire n4551;
  wire n4553;
  wire [3:0] n4555;
  wire n4557;
  wire [31:0] n4558;
  wire n4560;
  wire n4561;
  wire n4563;
  wire [3:0] n4565;
  wire n4567;
  wire [31:0] n4568;
  wire n4570;
  wire n4571;
  wire n4573;
  wire [3:0] n4575;
  wire n4577;
  wire [31:0] n4578;
  wire n4580;
  wire n4581;
  wire n4583;
  wire [3:0] n4585;
  wire [2:0] n4586;
  reg n4587;
  reg [3:0] n4588;
  wire n4590;
  wire [7:0] n4591;
  wire [7:0] n4592;
  wire n4602;
  wire n4604;
  wire [31:0] n4605;
  wire [31:0] n4607;
  wire [5:0] n4608;
  wire n4610;
  wire [31:0] n4611;
  wire [31:0] n4613;
  wire [5:0] n4614;
  wire n4616;
  wire [31:0] n4617;
  wire [31:0] n4619;
  wire [5:0] n4620;
  wire n4622;
  wire [31:0] n4623;
  wire [31:0] n4625;
  wire [5:0] n4626;
  wire n4628;
  wire [5:0] n4629;
  reg n4632;
  reg n4634;
  wire [79:0] n4635;
  reg [79:0] n4636;
  wire [79:0] n4637;
  reg [79:0] n4638;
  wire [79:0] n4639;
  reg [79:0] n4640;
  wire [79:0] n4641;
  reg [79:0] n4642;
  wire [79:0] n4643;
  reg [79:0] n4644;
  wire [79:0] n4645;
  reg [79:0] n4646;
  wire [79:0] n4647;
  reg [79:0] n4648;
  wire [79:0] n4649;
  reg [79:0] n4650;
  reg [31:0] n4652;
  reg [31:0] n4654;
  reg [31:0] n4656;
  reg [3:0] n4660;
  reg n4662;
  reg [5:0] n4663;
  reg [7:0] n4665;
  wire n4667;
  wire [31:0] n4668;
  wire [31:0] n4670;
  wire [5:0] n4671;
  wire n4673;
  wire [1:0] n4679;
  wire n4681;
  wire n4685;
  wire n4691;
  wire [15:0] n4692;
  wire n4694;
  wire [5:0] n4695;
  wire n4697;
  wire n4698;
  wire n4701;
  wire n4704;
  wire n4705;
  wire n4707;
  wire n4708;
  wire n4710;
  wire n4716;
  wire [1:0] n4724;
  wire n4726;
  wire [1:0] n4728;
  wire [1:0] n4729;
  wire [7:0] n4733;
  wire [31:0] n4735;
  wire [1:0] n4743;
  wire n4745;
  wire [1:0] n4747;
  wire [1:0] n4748;
  wire [7:0] n4752;
  wire [31:0] n4754;
  wire [1:0] n4755;
  wire n4757;
  wire n4760;
  wire [1:0] n4761;
  wire n4763;
  wire n4766;
  wire [31:0] n4767;
  wire n4772;
  wire n4774;
  wire [31:0] n4775;
  wire [31:0] n4777;
  wire [5:0] n4778;
  wire n4780;
  wire n4789;
  wire [31:0] n4790;
  wire [31:0] n4792;
  wire [5:0] n4793;
  wire n4795;
  wire n4797;
  wire n4798;
  wire [31:0] n4799;
  wire [31:0] n4801;
  wire [5:0] n4802;
  wire n4804;
  wire [31:0] n4805;
  wire [31:0] n4807;
  wire [5:0] n4808;
  wire n4810;
  wire [3:0] n4811;
  reg n4814;
  reg [3:0] n4817;
  reg [5:0] n4818;
  wire n4820;
  wire n4822;
  wire n4824;
  wire n4825;
  wire [31:0] n4826;
  wire n4828;
  wire [31:0] n4829;
  wire [31:0] n4831;
  wire [5:0] n4832;
  wire n4834;
  wire [3:0] n4836;
  wire [5:0] n4837;
  wire [31:0] n4838;
  wire [31:0] n4840;
  wire [5:0] n4841;
  wire n4842;
  wire n4843;
  wire [5:0] n4844;
  wire n4847;
  wire n4848;
  wire n4849;
  wire [31:0] n4850;
  wire [31:0] n4852;
  wire [5:0] n4853;
  wire n4856;
  wire n4857;
  wire n4858;
  wire [31:0] n4859;
  wire n4861;
  wire [31:0] n4862;
  wire [31:0] n4864;
  wire [5:0] n4865;
  wire n4867;
  wire [3:0] n4869;
  wire [5:0] n4870;
  wire n4872;
  wire [31:0] n4873;
  wire [31:0] n4875;
  wire [2:0] n4876;
  wire [2:0] n4878;
  wire [31:0] n4881;
  wire [31:0] n4883;
  wire [5:0] n4884;
  wire n4887;
  wire n4888;
  wire n4889;
  wire [31:0] n4890;
  wire [31:0] n4892;
  wire [2:0] n4893;
  wire [2:0] n4895;
  wire [31:0] n4898;
  wire [31:0] n4900;
  wire [5:0] n4901;
  wire n4904;
  wire n4905;
  wire n4906;
  wire [31:0] n4907;
  wire [31:0] n4909;
  wire [2:0] n4910;
  wire [2:0] n4912;
  wire [15:0] n4914;
  wire [31:0] n4916;
  wire [31:0] n4918;
  wire [30:0] n4919;
  wire [2:0] n4920;
  wire [31:0] n4921;
  wire [31:0] n4923;
  wire [2:0] n4924;
  wire [2:0] n4926;
  wire [63:0] n4928;
  wire [15:0] n4929;
  wire [79:0] n4930;
  wire [31:0] n4943;
  wire [31:0] n4945;
  wire [5:0] n4946;
  wire n4949;
  wire n4950;
  wire n4951;
  wire [31:0] n4952;
  wire n4954;
  wire [31:0] n4955;
  wire [31:0] n4957;
  wire [5:0] n4958;
  wire n4960;
  wire [3:0] n4962;
  wire [5:0] n4963;
  wire [2:0] n4964;
  reg n4965;
  reg n4970;
  reg [2:0] n4971;
  reg [79:0] n4972;
  reg n4975;
  reg [3:0] n4976;
  reg [5:0] n4977;
  reg [639:0] n4978;
  wire n4980;
  wire [31:0] n4981;
  wire n4983;
  wire [31:0] n4984;
  wire [31:0] n4986;
  wire [5:0] n4987;
  wire n4989;
  wire [3:0] n4991;
  wire [5:0] n4992;
  wire [1:0] n4993;
  reg n4994;
  reg n4998;
  reg [2:0] n4999;
  reg [79:0] n5000;
  reg n5002;
  reg [3:0] n5003;
  reg [5:0] n5004;
  reg [639:0] n5005;
  wire n5008;
  wire n5009;
  wire n5010;
  wire [6:0] n5011;
  reg n5013;
  reg n5014;
  wire [79:0] n5015;
  reg [79:0] n5016;
  wire [79:0] n5017;
  reg [79:0] n5018;
  wire [79:0] n5019;
  reg [79:0] n5020;
  wire [79:0] n5021;
  reg [79:0] n5022;
  wire [79:0] n5023;
  reg [79:0] n5024;
  wire [79:0] n5025;
  reg [79:0] n5026;
  wire [79:0] n5027;
  reg [79:0] n5028;
  wire [79:0] n5029;
  reg [79:0] n5030;
  reg n5034;
  reg [2:0] n5035;
  reg [79:0] n5036;
  reg n5038;
  reg [31:0] n5039;
  reg [31:0] n5041;
  reg [31:0] n5044;
  reg n5045;
  reg n5046;
  reg [3:0] n5050;
  reg n5051;
  reg [5:0] n5052;
  reg [7:0] n5053;
  reg [639:0] n5054;
  reg [7:0] n5055;
  wire n5056;
  wire n5057;
  wire [639:0] n5058;
  wire [639:0] n5059;
  wire n5063;
  wire [2:0] n5065;
  wire [79:0] n5066;
  wire n5068;
  wire [31:0] n5070;
  wire [31:0] n5072;
  wire [31:0] n5074;
  wire n5075;
  wire n5076;
  wire [3:0] n5078;
  wire n5079;
  wire [5:0] n5080;
  wire [7:0] n5081;
  wire [639:0] n5082;
  wire [7:0] n5083;
  wire n5085;
  wire n5088;
  wire n5091;
  wire n5094;
  wire n5097;
  wire n5100;
  wire n5103;
  wire n5106;
  wire n5109;
  wire [7:0] n5110;
  reg n5144;
  reg [2:0] n5153;
  reg [79:0] n5154;
  reg n5163;
  wire n5167;
  wire [2:0] n5168;
  wire [79:0] n5169;
  wire n5170;
  wire n5171;
  wire n5172;
  wire n5174;
  wire [3:0] n5176;
  wire n5178;
  wire n5180;
  wire n5182;
  wire n5184;
  wire [2:0] n5185;
  reg [31:0] n5187;
  wire [31:0] n5188;
  wire [1:0] n5194;
  wire n5196;
  wire n5200;
  wire n5206;
  wire [15:0] n5207;
  wire n5209;
  wire [5:0] n5210;
  wire n5212;
  wire n5213;
  wire n5216;
  wire n5219;
  wire n5220;
  wire n5222;
  wire n5223;
  wire n5225;
  wire n5231;
  wire [1:0] n5239;
  wire n5241;
  wire [1:0] n5243;
  wire [1:0] n5244;
  wire [7:0] n5248;
  wire [31:0] n5250;
  wire [1:0] n5258;
  wire n5260;
  wire [1:0] n5262;
  wire [1:0] n5263;
  wire [7:0] n5267;
  wire [31:0] n5269;
  wire [1:0] n5270;
  wire n5272;
  wire n5275;
  wire [1:0] n5276;
  wire n5278;
  wire n5281;
  wire [31:0] n5282;
  wire n5287;
  wire n5289;
  wire n5291;
  wire n5300;
  wire n5302;
  wire [2:0] n5303;
  reg [31:0] n5304;
  reg [31:0] n5306;
  reg [31:0] n5309;
  reg n5312;
  reg n5313;
  wire [31:0] n5316;
  wire [31:0] n5318;
  wire [31:0] n5320;
  wire n5322;
  wire n5323;
  wire n5325;
  wire n5326;
  wire n5328;
  wire [3:0] n5330;
  wire n5332;
  wire [12:0] n5333;
  reg [31:0] n5337;
  reg n5342;
  reg n5344;
  reg [639:0] n5346;
  reg n5352;
  reg [2:0] n5354;
  reg [79:0] n5356;
  reg n5360;
  wire [5:0] n5361;
  wire [5:0] n5362;
  wire [5:0] n5363;
  wire [5:0] n5364;
  reg [5:0] n5366;
  wire [1:0] n5367;
  wire [1:0] n5368;
  wire [1:0] n5369;
  wire [1:0] n5370;
  reg [1:0] n5372;
  wire [5:0] n5373;
  wire [5:0] n5374;
  wire [5:0] n5375;
  wire [5:0] n5376;
  reg [5:0] n5378;
  wire [1:0] n5379;
  wire [1:0] n5380;
  wire [1:0] n5381;
  wire [1:0] n5382;
  reg [1:0] n5384;
  wire [15:0] n5385;
  wire [15:0] n5386;
  wire [15:0] n5387;
  wire [15:0] n5388;
  reg [15:0] n5390;
  wire [12:0] n5395;
  wire [12:0] n5396;
  wire [12:0] n5397;
  wire [12:0] n5398;
  wire [12:0] n5399;
  reg [12:0] n5401;
  wire n5402;
  wire n5403;
  wire n5404;
  wire n5405;
  wire n5406;
  reg n5408;
  wire n5409;
  wire n5410;
  wire n5411;
  wire n5412;
  wire n5413;
  wire n5414;
  reg n5416;
  wire n5417;
  wire n5418;
  wire n5419;
  wire n5420;
  wire n5421;
  wire n5422;
  reg n5424;
  wire n5425;
  wire n5426;
  wire n5427;
  wire n5428;
  wire n5429;
  wire n5430;
  reg n5432;
  wire n5433;
  wire n5434;
  wire n5435;
  wire n5436;
  wire n5437;
  wire n5438;
  reg n5440;
  wire n5441;
  wire n5442;
  wire n5443;
  wire n5444;
  wire n5445;
  wire n5446;
  reg n5448;
  wire [1:0] n5449;
  wire [1:0] n5450;
  wire [1:0] n5451;
  wire [1:0] n5452;
  wire [1:0] n5453;
  wire [1:0] n5454;
  reg [1:0] n5456;
  wire n5457;
  wire n5458;
  wire n5459;
  wire n5460;
  wire n5461;
  wire n5462;
  reg n5464;
  wire n5465;
  wire n5466;
  wire n5467;
  wire n5468;
  wire n5469;
  wire n5470;
  reg n5472;
  wire n5473;
  wire n5474;
  wire n5475;
  wire n5476;
  wire n5477;
  wire n5478;
  reg n5480;
  wire n5481;
  wire n5482;
  wire n5483;
  wire n5484;
  wire n5485;
  wire n5486;
  reg n5488;
  wire n5489;
  wire n5490;
  wire n5491;
  wire n5492;
  wire n5493;
  wire n5494;
  reg n5496;
  wire n5497;
  wire n5498;
  wire n5499;
  wire n5500;
  wire n5501;
  wire n5502;
  reg n5504;
  wire n5505;
  wire n5506;
  wire n5507;
  wire n5508;
  wire n5509;
  reg n5511;
  wire [3:0] n5512;
  wire [3:0] n5513;
  wire [3:0] n5514;
  wire [3:0] n5515;
  wire [3:0] n5516;
  reg [3:0] n5518;
  reg [31:0] n5522;
  reg n5526;
  reg n5528;
  reg [1:0] n5530;
  reg n5534;
  reg [15:0] n5536;
  reg [31:0] n5538;
  reg [3:0] n5544;
  reg [7:0] n5548;
  reg n5551;
  reg [7:0] n5553;
  reg n5555;
  reg [7:0] n5559;
  reg [5:0] n5561;
  reg [7:0] n5563;
  reg [639:0] n5569;
  reg [7:0] n5571;
  reg n5574;
  reg [6:0] n5576;
  reg [79:0] n5578;
  reg [79:0] n5580;
  reg n5583;
  reg [6:0] n5585;
  reg [79:0] n5587;
  reg [79:0] n5589;
  reg n5591;
  reg n5593;
  reg n5595;
  reg n5597;
  reg [79:0] n5599;
  reg n5601;
  reg [2:0] n5603;
  reg [2:0] n5605;
  reg [95:0] n5607;
  reg [6:0] n5609;
  reg n5611;
  reg n5613;
  reg n5615;
  reg [5:0] n5623;
  reg [31:0] n5625;
  wire n5626;
  wire [30:0] n5627;
  wire [31:0] n5628;
  wire n5630;
  wire n5631;
  wire n5633;
  wire [7:0] n5635;
  wire n5637;
  wire n5639;
  wire n5641;
  wire n5643;
  wire n5645;
  wire n5647;
  wire n5648;
  wire [4:0] n5649;
  reg n5655;
  reg [7:0] n5661;
  wire n5662;
  wire [7:0] n5663;
  wire [31:0] n5664;
  wire n5666;
  wire [7:0] n5669;
  wire [7:0] n5671;
  wire n5673;
  wire [7:0] n5674;
  wire [31:0] n5675;
  wire n5677;
  wire n5679;
  wire [7:0] n5681;
  wire n5683;
  wire n5685;
  wire n5687;
  wire n5689;
  wire [3:0] n5691;
  wire n5693;
  wire n5695;
  wire n5697;
  wire [3:0] n5699;
  wire [31:0] n5711;
  wire [31:0] n5715;
  wire n5934;
  wire n5937;
  wire [2:0] n5940;
  wire [79:0] n5944;
  wire n5953;
  wire n5956;
  reg n5959;
  wire n5967;
  wire [2:0] n5971;
  wire n5980;
  wire n5981;
  wire n5982;
  wire n5983;
  wire n5987;
  wire n5991;
  wire n5992;
  wire [31:0] n5993;
  wire [31:0] n5995;
  wire [9:0] n5996;
  wire [31:0] n5997;
  wire n5999;
  wire n6005;
  wire [9:0] n6007;
  wire n6010;
  wire [9:0] n6012;
  wire n6013;
  wire n6014;
  wire n6026;
  wire n6048;
  wire n6081;
  wire [2:0] n6082;
  reg [15:0] n6083;
  reg n6087;
  wire n6096;
  wire n6103;
  wire n6105;
  wire n6107;
  wire n6108;
  wire n6109;
  wire n6110;
  wire n6112;
  wire n6113;
  wire [2:0] n6115;
  wire n6117;
  wire [31:0] n6118;
  wire [31:0] n6120;
  wire [9:0] n6121;
  wire [30:0] n6122;
  wire [31:0] n6123;
  wire n6125;
  wire n6127;
  wire n6129;
  wire n6130;
  wire n6131;
  wire n6132;
  wire n6134;
  wire n6136;
  wire n6137;
  wire n6139;
  wire n6140;
  wire n6141;
  wire [2:0] n6144;
  wire [2:0] n6148;
  wire [2:0] n6152;
  wire [31:0] n6155;
  wire n6157;
  wire [2:0] n6159;
  wire n6163;
  wire [31:0] n6164;
  wire [31:0] n6166;
  wire [9:0] n6167;
  wire [2:0] n6185;
  wire [2:0] n6191;
  wire [31:0] n6196;
  wire n6198;
  wire [2:0] n6200;
  wire n6204;
  wire n6206;
  wire n6207;
  wire n6208;
  wire n6209;
  wire [2:0] n6211;
  wire [31:0] n6212;
  wire n6214;
  wire [2:0] n6216;
  wire n6220;
  wire n6222;
  wire [31:0] n6223;
  wire n6225;
  wire [31:0] n6226;
  wire [31:0] n6228;
  wire [9:0] n6229;
  wire [9:0] n6230;
  wire [2:0] n6232;
  wire n6238;
  wire [6:0] n6239;
  reg [9:0] n6242;
  reg [2:0] n6250;
  wire n6263;
  wire n6265;
  wire n6267;
  wire n6269;
  wire n6270;
  reg [15:0] n6273;
  wire n6275;
  wire n6277;
  wire [1:0] n6278;
  reg [15:0] n6281;
  wire n6283;
  wire n6285;
  wire n6287;
  wire n6289;
  wire [15:0] n6292;
  wire [15:0] n6294;
  wire [15:0] n6296;
  wire [15:0] n6298;
  wire [15:0] n6299;
  wire n6301;
  wire n6303;
  wire n6304;
  wire n6305;
  wire [31:0] n6306;
  wire n6308;
  wire [15:0] n6311;
  wire [15:0] n6313;
  wire n6315;
  wire n6317;
  wire n6319;
  wire n6321;
  wire n6322;
  wire n6323;
  wire [31:0] n6324;
  wire n6326;
  wire [15:0] n6329;
  wire [15:0] n6331;
  wire [15:0] n6333;
  wire n6335;
  wire n6337;
  wire n6339;
  wire [6:0] n6343;
  reg [15:0] n6349;
  wire n6350;
  localparam [15:0] n6351 = 16'b0000000000000000;
  wire [11:0] n6352;
  wire n6354;
  wire n6356;
  wire n6358;
  wire n6360;
  wire n6362;
  wire n6363;
  wire n6365;
  wire n6366;
  wire n6367;
  wire n6369;
  wire n6371;
  wire n6373;
  wire [2:0] n6374;
  reg [15:0] n6379;
  wire [15:0] n6381;
  wire n6384;
  wire [15:0] n6385;
  wire n6530;
  wire n6532;
  wire n6534;
  wire n6536;
  wire n6538;
  wire n6540;
  wire n6542;
  wire [15:0] n6543;
  wire n6545;
  wire [15:0] n6546;
  wire n6548;
  wire [8:0] n6549;
  reg [15:0] n6554;
  wire n6556;
  reg n6557;
  wire n6558;
  wire n6559;
  wire n6560;
  reg n6561;
  wire n6562;
  reg n6563;
  wire [639:0] n6564;
  reg [639:0] n6565;
  wire n6570;
  reg n6571;
  wire [2:0] n6572;
  reg [2:0] n6573;
  wire [79:0] n6574;
  reg [79:0] n6575;
  wire n6582;
  reg n6583;
  wire [31:0] n6588;
  reg [31:0] n6589;
  wire [31:0] n6594;
  reg [31:0] n6595;
  wire [31:0] n6598;
  reg [31:0] n6599;
  wire n6602;
  wire n6603;
  wire n6604;
  reg n6605;
  wire n6606;
  wire n6607;
  wire n6608;
  reg n6609;
  wire n6610;
  wire n6611;
  wire [1:0] n6612;
  reg [1:0] n6613;
  wire [15:0] n6618;
  reg [15:0] n6619;
  wire [15:0] n6620;
  reg [15:0] n6621;
  wire [15:0] n6622;
  reg [15:0] n6623;
  wire [15:0] n6624;
  reg [15:0] n6625;
  wire n6630;
  reg n6631;
  wire n6632;
  reg n6633;
  wire n6634;
  reg n6635;
  wire [9:0] n6636;
  reg [9:0] n6637;
  reg [9:0] n6638;
  wire n6639;
  reg n6640;
  wire n6643;
  wire n6644;
  wire n6645;
  reg n6646;
  wire n6653;
  wire n6654;
  wire n6655;
  reg n6656;
  wire [2:0] n6657;
  reg [2:0] n6658;
  wire n6661;
  wire n6662;
  wire [2:0] n6663;
  reg [2:0] n6664;
  wire n6677;
  wire n6678;
  wire [15:0] n6679;
  reg [15:0] n6680;
  wire n6681;
  wire n6682;
  wire [31:0] n6683;
  reg [31:0] n6684;
  wire [3:0] n6685;
  reg [3:0] n6686;
  wire n6687;
  reg n6688;
  wire [7:0] n6691;
  reg [7:0] n6692;
  wire n6693;
  reg n6694;
  wire [7:0] n6695;
  reg [7:0] n6696;
  wire n6697;
  reg n6698;
  wire [7:0] n6699;
  reg [7:0] n6700;
  wire [5:0] n6701;
  reg [5:0] n6702;
  wire [7:0] n6703;
  reg [7:0] n6704;
  wire n6709;
  wire n6710;
  wire [639:0] n6711;
  reg [639:0] n6712;
  wire [6:0] n6713;
  reg [6:0] n6714;
  wire [2:0] n6715;
  reg [2:0] n6716;
  wire [2:0] n6717;
  reg [2:0] n6718;
  wire [2:0] n6719;
  reg [2:0] n6720;
  wire [2:0] n6721;
  reg [2:0] n6722;
  wire [2:0] n6723;
  reg [2:0] n6724;
  wire [7:0] n6728;
  reg [7:0] n6729;
  wire n6730;
  wire n6731;
  wire n6732;
  reg n6733;
  wire n6734;
  wire n6735;
  wire [6:0] n6736;
  reg [6:0] n6737;
  wire n6738;
  wire n6739;
  wire [79:0] n6740;
  reg [79:0] n6741;
  wire n6742;
  wire n6743;
  wire [79:0] n6744;
  reg [79:0] n6745;
  wire n6746;
  wire n6747;
  wire n6748;
  reg n6749;
  wire n6750;
  wire n6751;
  wire [6:0] n6752;
  reg [6:0] n6753;
  wire n6754;
  wire n6755;
  wire [79:0] n6756;
  reg [79:0] n6757;
  wire n6758;
  wire n6759;
  wire [79:0] n6760;
  reg [79:0] n6761;
  wire n6762;
  wire n6763;
  wire n6764;
  reg n6765;
  wire n6766;
  wire n6767;
  wire n6768;
  reg n6769;
  wire n6770;
  wire n6771;
  wire n6772;
  reg n6773;
  wire n6774;
  wire n6775;
  wire n6776;
  reg n6777;
  wire n6778;
  wire n6779;
  wire [79:0] n6780;
  reg [79:0] n6781;
  wire n6783;
  wire n6784;
  wire n6785;
  reg n6786;
  wire n6787;
  wire n6788;
  wire [2:0] n6789;
  reg [2:0] n6790;
  wire n6791;
  wire n6792;
  wire [2:0] n6793;
  reg [2:0] n6794;
  wire n6795;
  wire n6796;
  wire [95:0] n6797;
  reg [95:0] n6798;
  wire n6799;
  wire n6800;
  wire [6:0] n6801;
  reg [6:0] n6802;
  wire n6803;
  wire n6804;
  wire n6805;
  reg n6806;
  reg n6807;
  wire n6808;
  reg n6809;
  wire n6810;
  reg n6811;
  wire n6812;
  wire n6813;
  wire [79:0] n6814;
  reg [79:0] n6815;
  wire n6832;
  wire n6833;
  wire [5:0] n6834;
  reg [5:0] n6835;
  wire n6836;
  wire n6837;
  wire [31:0] n6838;
  reg [31:0] n6839;
  wire [31:0] n6840;
  reg [31:0] n6841;
  wire n6842;
  wire n6843;
  wire n6844;
  wire n6845;
  wire n6846;
  wire n6847;
  wire n6848;
  wire n6849;
  wire n6850;
  wire n6851;
  wire n6852;
  wire n6853;
  wire n6854;
  wire n6855;
  wire n6856;
  wire n6857;
  wire n6858;
  wire n6859;
  wire [79:0] n6860;
  wire [79:0] n6861;
  wire [79:0] n6862;
  wire [79:0] n6863;
  wire [79:0] n6864;
  wire [79:0] n6865;
  wire [79:0] n6866;
  wire [79:0] n6867;
  wire [79:0] n6868;
  wire [79:0] n6869;
  wire [79:0] n6870;
  wire [79:0] n6871;
  wire [79:0] n6872;
  wire [79:0] n6873;
  wire [79:0] n6874;
  wire [79:0] n6875;
  wire [639:0] n6876;
  wire [9:0] n6878;
  wire [9:0] n6879;
  wire [560:0] n6880;
  wire [639:0] n6882;
  wire [79:0] n6883;
  wire n6884;
  wire [9:0] n6886;
  wire [9:0] n6887;
  wire [79:0] n6888;
  wire [79:0] n6889;
  wire [560:0] n6890;
  wire [639:0] n6892;
  wire [79:0] n6893;
  wire n6894;
  wire [9:0] n6896;
  wire [9:0] n6897;
  wire [9:0] n6899;
  wire [9:0] n6900;
  wire [560:0] n6901;
  wire [639:0] n6903;
  wire [79:0] n6904;
  wire n6905;
  wire [574:0] n6906;
  wire [639:0] n6908;
  wire [79:0] n6909;
  wire [9:0] n6910;
  wire [595:0] n6911;
  wire [639:0] n6913;
  wire [79:0] n6914;
  wire [19:0] n6915;
  wire [9:0] n6917;
  wire [9:0] n6918;
  wire [9:0] n6920;
  wire [9:0] n6921;
  wire [560:0] n6922;
  wire [639:0] n6924;
  wire [79:0] n6925;
  wire n6926;
  wire [9:0] n6928;
  wire [9:0] n6929;
  wire [9:0] n6931;
  wire [9:0] n6932;
  wire [560:0] n6933;
  wire [639:0] n6935;
  wire [79:0] n6936;
  wire n6937;
  wire [9:0] n6939;
  wire [9:0] n6940;
  wire [9:0] n6942;
  wire [9:0] n6943;
  wire [9:0] n6945;
  wire [9:0] n6946;
  wire [9:0] n6948;
  wire [9:0] n6949;
  wire [9:0] n6951;
  wire [9:0] n6952;
  wire [560:0] n6953;
  wire [639:0] n6955;
  wire [79:0] n6956;
  wire n6957;
  wire [79:0] n6958;
  wire [79:0] n6959;
  wire [79:0] n6960;
  wire [9:0] n6962;
  wire [9:0] n6963;
  wire [9:0] n6965;
  wire [9:0] n6966;
  wire [79:0] n6967;
  wire [15:0] n6968;
  wire n6969;
  wire n6970;
  wire n6971;
  wire n6972;
  wire n6973;
  wire n6974;
  wire n6975;
  wire n6976;
  wire n6977;
  wire n6978;
  wire n6979;
  wire n6980;
  wire n6981;
  wire n6982;
  wire n6983;
  wire n6984;
  wire n6985;
  wire n6986;
  wire [47:0] n6987;
  wire [31:0] n6988;
  wire [31:0] n6989;
  wire [47:0] n6990;
  wire [31:0] n6991;
  wire [31:0] n6992;
  wire [47:0] n6993;
  wire [31:0] n6994;
  wire [31:0] n6995;
  wire [47:0] n6996;
  wire [31:0] n6997;
  wire [31:0] n6998;
  wire [47:0] n6999;
  wire [31:0] n7000;
  wire [31:0] n7001;
  wire [47:0] n7002;
  wire [31:0] n7003;
  wire [31:0] n7004;
  wire [47:0] n7005;
  wire [31:0] n7006;
  wire [31:0] n7007;
  wire [47:0] n7008;
  wire [31:0] n7009;
  wire [31:0] n7010;
  wire [639:0] n7011;
  wire n7012;
  wire n7013;
  wire n7014;
  wire n7015;
  wire n7016;
  wire n7017;
  wire n7018;
  wire n7019;
  wire n7020;
  wire n7021;
  wire n7022;
  wire n7023;
  wire n7024;
  wire n7025;
  wire n7026;
  wire n7027;
  wire n7028;
  wire n7029;
  wire [15:0] n7030;
  wire [31:0] n7031;
  wire [31:0] n7032;
  wire [47:0] n7033;
  wire [31:0] n7034;
  wire [31:0] n7035;
  wire [47:0] n7036;
  wire [31:0] n7037;
  wire [31:0] n7038;
  wire [47:0] n7039;
  wire [31:0] n7040;
  wire [31:0] n7041;
  wire [47:0] n7042;
  wire [31:0] n7043;
  wire [31:0] n7044;
  wire [47:0] n7045;
  wire [31:0] n7046;
  wire [31:0] n7047;
  wire [47:0] n7048;
  wire [31:0] n7049;
  wire [31:0] n7050;
  wire [47:0] n7051;
  wire [31:0] n7052;
  wire [31:0] n7053;
  wire [31:0] n7054;
  wire [639:0] n7055;
  wire n7056;
  wire n7057;
  wire n7058;
  wire n7059;
  wire n7060;
  wire n7061;
  wire n7062;
  wire n7063;
  wire n7064;
  wire n7065;
  wire n7066;
  wire n7067;
  wire n7068;
  wire n7069;
  wire n7070;
  wire n7071;
  wire n7072;
  wire n7073;
  wire [15:0] n7074;
  wire [15:0] n7075;
  wire [63:0] n7076;
  wire [15:0] n7077;
  wire [15:0] n7078;
  wire [63:0] n7079;
  wire [15:0] n7080;
  wire [15:0] n7081;
  wire [63:0] n7082;
  wire [15:0] n7083;
  wire [15:0] n7084;
  wire [63:0] n7085;
  wire [15:0] n7086;
  wire [15:0] n7087;
  wire [63:0] n7088;
  wire [15:0] n7089;
  wire [15:0] n7090;
  wire [63:0] n7091;
  wire [15:0] n7092;
  wire [15:0] n7093;
  wire [63:0] n7094;
  wire [15:0] n7095;
  wire [15:0] n7096;
  wire [63:0] n7097;
  wire [639:0] n7098;
  wire [9:0] n7100;
  wire [9:0] n7101;
  wire [79:0] n7102;
  assign fpu_data_out = n6841; //(module output)
  assign fmovem_data_out = \fpu_movem.fmovem_data_out ; //(module output)
  assign fpu_busy = fpu_busy_internal; //(module output)
  assign fpu_done = fpu_done_i; //(module output)
  assign fpu_exception = fpu_exception_i; //(module output)
  assign exception_code = n197; //(module output)
  assign fpcr_out = fpcr; //(module output)
  assign fpsr_out = n196; //(module output)
  assign fpiar_out = fpiar; //(module output)
  assign fsave_frame_size = fsave_frame_size_internal; //(module output)
  assign fsave_size_valid = fsave_size_valid_internal; //(module output)
  assign cir_data_out = n6554; //(module output)
  assign cir_data_valid = cir_data_valid_i; //(module output)
  /* TG68K_FPU.vhd:86:16  */
  always @*
    fpu_done_i = n6557; // (isignal)
  initial
    fpu_done_i = 1'b0;
  /* TG68K_FPU.vhd:87:16  */
  always @*
    fpu_exception_i = n6561; // (isignal)
  initial
    fpu_exception_i = 1'b0;
  /* TG68K_FPU.vhd:88:16  */
  always @*
    cir_data_valid_i = n6563; // (isignal)
  initial
    cir_data_valid_i = 1'b0;
  /* TG68K_FPU.vhd:97:16  */
  assign fp_registers = n6565; // (signal)
  /* TG68K_FPU.vhd:100:16  */
  always @*
    fp_reg_write_enable = n6571; // (isignal)
  initial
    fp_reg_write_enable = 1'b0;
  /* TG68K_FPU.vhd:101:16  */
  always @*
    fp_reg_write_addr = n6573; // (isignal)
  initial
    fp_reg_write_addr = 3'b000;
  /* TG68K_FPU.vhd:102:16  */
  always @*
    fp_reg_write_data = n6575; // (isignal)
  initial
    fp_reg_write_data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:105:16  */
  always @*
    fp_reg_access_valid = n6583; // (isignal)
  initial
    fp_reg_access_valid = 1'b0;
  /* TG68K_FPU.vhd:129:16  */
  always @*
    fpcr = n6589; // (isignal)
  initial
    fpcr = 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:138:16  */
  always @*
    fpsr = n6595; // (isignal)
  initial
    fpsr = 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:141:16  */
  always @*
    fpiar = n6599; // (isignal)
  initial
    fpiar = 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:143:16  */
  always @*
    fpcr_rounding_mode_valid = n6605; // (isignal)
  initial
    fpcr_rounding_mode_valid = 1'b1;
  /* TG68K_FPU.vhd:144:16  */
  always @*
    fpcr_precision_valid = n6609; // (isignal)
  initial
    fpcr_precision_valid = 1'b1;
  /* TG68K_FPU.vhd:145:16  */
  assign fpcr_precision_bits = n6613; // (signal)
  /* TG68K_FPU.vhd:154:16  */
  always @*
    response_cir = n6619; // (isignal)
  initial
    response_cir = 16'b0000000000000000;
  /* TG68K_FPU.vhd:155:16  */
  always @*
    command_cir = n6621; // (isignal)
  initial
    command_cir = 16'b0000000000000000;
  /* TG68K_FPU.vhd:156:16  */
  always @*
    condition_cir = n6623; // (isignal)
  initial
    condition_cir = 16'b0000000000000000;
  /* TG68K_FPU.vhd:157:16  */
  always @*
    save_cir = n6625; // (isignal)
  initial
    save_cir = 16'b0000000000000000;
  /* TG68K_FPU.vhd:160:16  */
  always @*
    cir_read_reg = n6631; // (isignal)
  initial
    cir_read_reg = 1'b0;
  /* TG68K_FPU.vhd:163:16  */
  always @*
    cir_write_reg = n6633; // (isignal)
  initial
    cir_write_reg = 1'b0;
  /* TG68K_FPU.vhd:164:16  */
  always @*
    cir_read_active = n6635; // (isignal)
  initial
    cir_read_active = 1'b0;
  /* TG68K_FPU.vhd:165:16  */
  always @*
    cir_timeout_counter = n6637; // (isignal)
  initial
    cir_timeout_counter = 10'b0000000000;
  /* TG68K_FPU.vhd:166:16  */
  always @*
    state_timeout_counter = n6638; // (isignal)
  initial
    state_timeout_counter = 10'b0000000000;
  /* TG68K_FPU.vhd:167:16  */
  always @*
    command_pending = n6640; // (isignal)
  initial
    command_pending = 1'b0;
  /* TG68K_FPU.vhd:168:16  */
  always @*
    command_valid = 1'b0; // (isignal)
  initial
    command_valid = 1'b0;
  /* TG68K_FPU.vhd:170:16  */
  always @*
    restore_privilege_violation = n6646; // (isignal)
  initial
    restore_privilege_violation = 1'b0;
  /* TG68K_FPU.vhd:174:16  */
  always @*
    cir_address_error = n6656; // (isignal)
  initial
    cir_address_error = 1'b0;
  /* TG68K_FPU.vhd:175:16  */
  always @*
    current_privilege_level = n6658; // (isignal)
  initial
    current_privilege_level = 3'b000;
  /* TG68K_FPU.vhd:178:16  */
  always @*
    cir_handshake_state = n6664; // (isignal)
  initial
    cir_handshake_state = 3'b000;
  /* TG68K_FPU.vhd:184:16  */
  always @*
    operation_word_cir = n6680; // (isignal)
  initial
    operation_word_cir = 16'b0000000000000000;
  /* TG68K_FPU.vhd:185:16  */
  always @*
    command_address_cir = n6684; // (isignal)
  initial
    command_address_cir = 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:203:16  */
  always @*
    fpu_state = n6686; // (isignal)
  initial
    fpu_state = 4'b0000;
  /* TG68K_FPU.vhd:205:16  */
  always @*
    fpu_busy_internal = n6688; // (isignal)
  initial
    fpu_busy_internal = 1'b0;
  /* TG68K_FPU.vhd:208:16  */
  assign fsave_frame_format = n285; // (signal)
  /* TG68K_FPU.vhd:211:16  */
  always @*
    fsave_frame_size_internal = n287; // (isignal)
  initial
    fsave_frame_size_internal = 8'b00111100;
  /* TG68K_FPU.vhd:212:16  */
  always @*
    fsave_size_valid_internal = 1'b1; // (isignal)
  initial
    fsave_size_valid_internal = 1'b1;
  /* TG68K_FPU.vhd:214:16  */
  always @*
    fsave_frame_format_latched = n6692; // (isignal)
  initial
    fsave_frame_format_latched = 8'b01100000;
  /* TG68K_FPU.vhd:216:16  */
  always @*
    fpu_just_reset = n6694; // (isignal)
  initial
    fpu_just_reset = 1'b0;
  /* TG68K_FPU.vhd:219:16  */
  assign movem_register_list = n6696; // (signal)
  /* TG68K_FPU.vhd:220:16  */
  assign movem_direction = n6698; // (signal)
  /* TG68K_FPU.vhd:223:16  */
  always @*
    timeout_counter = n6700; // (isignal)
  initial
    timeout_counter = 8'b00000000;
  /* TG68K_FPU.vhd:246:16  */
  always @*
    fsave_counter = n6702; // (isignal)
  initial
    fsave_counter = 6'b000000;
  /* TG68K_FPU.vhd:247:16  */
  assign frestore_frame_format = n6704; // (signal)
  /* TG68K_FPU.vhd:254:16  */
  assign frestore_fp_temp = n6712; // (signal)
  /* TG68K_FPU.vhd:257:16  */
  assign decoder_instruction_type = fpu_decoder_n81; // (signal)
  /* TG68K_FPU.vhd:258:16  */
  assign decoder_operation_code = fpu_decoder_n82; // (signal)
  /* TG68K_FPU.vhd:259:16  */
  assign decoder_source_format = fpu_decoder_n83; // (signal)
  /* TG68K_FPU.vhd:260:16  */
  assign decoder_dest_format = fpu_decoder_n84; // (signal)
  /* TG68K_FPU.vhd:261:16  */
  assign decoder_source_reg = fpu_decoder_n85; // (signal)
  /* TG68K_FPU.vhd:262:16  */
  assign decoder_dest_reg = fpu_decoder_n86; // (signal)
  /* TG68K_FPU.vhd:263:16  */
  assign decoder_ea_mode = fpu_decoder_n87; // (signal)
  /* TG68K_FPU.vhd:264:16  */
  assign decoder_ea_register = fpu_decoder_n88; // (signal)
  /* TG68K_FPU.vhd:266:16  */
  assign decoder_valid_instruction = fpu_decoder_n90; // (signal)
  /* TG68K_FPU.vhd:268:16  */
  assign decoder_illegal = fpu_decoder_n92; // (signal)
  /* TG68K_FPU.vhd:269:16  */
  assign decoder_unsupported = fpu_decoder_n93; // (signal)
  /* TG68K_FPU.vhd:272:16  */
  assign fpu_operation = n6714; // (signal)
  /* TG68K_FPU.vhd:273:16  */
  assign source_reg = n6716; // (signal)
  /* TG68K_FPU.vhd:274:16  */
  assign dest_reg = n6718; // (signal)
  /* TG68K_FPU.vhd:275:16  */
  assign data_format = n6720; // (signal)
  /* TG68K_FPU.vhd:276:16  */
  assign ea_mode = n6722; // (signal)
  /* TG68K_FPU.vhd:277:16  */
  assign ea_register = n6724; // (signal)
  /* TG68K_FPU.vhd:283:16  */
  assign exception_code_internal = n6729; // (signal)
  /* TG68K_FPU.vhd:286:16  */
  assign alu_start_operation = n6733; // (signal)
  /* TG68K_FPU.vhd:287:16  */
  assign alu_operation_code = n6737; // (signal)
  /* TG68K_FPU.vhd:288:16  */
  assign alu_operand_a = n6741; // (signal)
  /* TG68K_FPU.vhd:289:16  */
  assign alu_operand_b = n6745; // (signal)
  /* TG68K_FPU.vhd:300:16  */
  assign exception_reset = n190; // (signal)
  /* TG68K_FPU.vhd:301:16  */
  assign exception_op_valid = n191; // (signal)
  /* TG68K_FPU.vhd:302:16  */
  assign exception_op_type = n193; // (signal)
  /* TG68K_FPU.vhd:310:16  */
  assign trans_start_operation = n6749; // (signal)
  /* TG68K_FPU.vhd:311:16  */
  assign trans_operation_code = n6753; // (signal)
  /* TG68K_FPU.vhd:312:16  */
  assign trans_operand = n6757; // (signal)
  /* TG68K_FPU.vhd:313:16  */
  assign trans_result = fpu_trans_n129; // (signal)
  /* TG68K_FPU.vhd:314:16  */
  assign trans_result_valid = fpu_trans_n130; // (signal)
  /* TG68K_FPU.vhd:315:16  */
  assign trans_overflow = fpu_trans_n131; // (signal)
  /* TG68K_FPU.vhd:316:16  */
  assign trans_underflow = fpu_trans_n132; // (signal)
  /* TG68K_FPU.vhd:317:16  */
  assign trans_inexact = fpu_trans_n133; // (signal)
  /* TG68K_FPU.vhd:318:16  */
  assign trans_invalid = fpu_trans_n134; // (signal)
  /* TG68K_FPU.vhd:320:16  */
  assign trans_operation_done = fpu_trans_n136; // (signal)
  /* TG68K_FPU.vhd:324:16  */
  assign final_result = n6761; // (signal)
  /* TG68K_FPU.vhd:325:16  */
  assign final_overflow = n6765; // (signal)
  /* TG68K_FPU.vhd:326:16  */
  assign final_underflow = n6769; // (signal)
  /* TG68K_FPU.vhd:327:16  */
  assign final_inexact = n6773; // (signal)
  /* TG68K_FPU.vhd:328:16  */
  assign final_invalid = n6777; // (signal)
  /* TG68K_FPU.vhd:333:16  */
  assign result_data = n6781; // (signal)
  /* TG68K_FPU.vhd:337:16  */
  assign converter_start = n6786; // (signal)
  /* TG68K_FPU.vhd:340:16  */
  assign converter_source_format = n6790; // (signal)
  /* TG68K_FPU.vhd:341:16  */
  assign converter_dest_format = n6794; // (signal)
  /* TG68K_FPU.vhd:342:16  */
  assign converter_data_in = n6798; // (signal)
  /* TG68K_FPU.vhd:350:16  */
  assign rom_offset = n6802; // (signal)
  /* TG68K_FPU.vhd:351:16  */
  assign rom_read_enable = n6806; // (signal)
  /* TG68K_FPU.vhd:352:16  */
  assign constrom_result = fpu_const_rom_n173; // (signal)
  /* TG68K_FPU.vhd:353:16  */
  assign constrom_valid = fpu_const_rom_n174; // (signal)
  /* TG68K_FPU.vhd:356:16  */
  assign movem_start = n6807; // (signal)
  /* TG68K_FPU.vhd:359:16  */
  always @*
    movem_predecrement = n6809; // (isignal)
  initial
    movem_predecrement = 1'b0;
  /* TG68K_FPU.vhd:360:16  */
  always @*
    movem_postincrement = n6811; // (isignal)
  initial
    movem_postincrement = 1'b0;
  /* TG68K_FPU.vhd:375:16  */
  assign movem_reg_data_in = n6815; // (signal)
  /* TG68K_FPU.vhd:386:16  */
  assign fp_to_int_shift = n6835; // (signal)
  /* TG68K_FPU.vhd:387:16  */
  assign fp_to_int_result = n6839; // (signal)
  /* TG68K_FPU.vhd:750:9  */
  tg68k_fpu_decoder fpu_decoder (
    .clk(clk),
    .nreset(nReset),
    .opcode(opcode),
    .extension_word(extension_word),
    .decode_enable(fpu_enable),
    .instruction_type(fpu_decoder_n81),
    .operation_code(fpu_decoder_n82),
    .source_format(fpu_decoder_n83),
    .dest_format(fpu_decoder_n84),
    .source_reg(fpu_decoder_n85),
    .dest_reg(fpu_decoder_n86),
    .ea_mode(fpu_decoder_n87),
    .ea_register(fpu_decoder_n88),
    .needs_extension_word(),
    .valid_instruction(fpu_decoder_n90),
    .privileged_instruction(),
    .illegal_instruction(fpu_decoder_n92),
    .unsupported_instruction(fpu_decoder_n93));
  /* TG68K_FPU.vhd:784:9  */
  tg68k_fpu_alu fpu_alu (
    .clk(clk),
    .nreset(nReset),
    .clkena(clkena),
    .start_operation(alu_start_operation),
    .operation_code(alu_operation_code),
    .rounding_mode(n118),
    .operand_a(alu_operand_a),
    .operand_b(alu_operand_b),
    .result(alu_result),
    .result_valid(alu_result_valid),
    .overflow(alu_overflow),
    .underflow(alu_underflow),
    .inexact(alu_inexact),
    .invalid(alu_invalid),
    .divide_by_zero(alu_divide_by_zero),
    .quotient_byte(alu_quotient_byte),
    .operation_busy(),
    .operation_done(alu_operation_done));
  /* TG68K_FPU.vhd:793:38  */
  assign n118 = fpcr[15:14]; // extract
  /* TG68K_FPU.vhd:819:9  */
  tg68k_fpu_transcendental fpu_trans (
    .clk(clk),
    .nreset(nReset),
    .clkena(clkena),
    .start_operation(trans_start_operation),
    .operation_code(trans_operation_code),
    .operand(trans_operand),
    .result(fpu_trans_n129),
    .result_valid(fpu_trans_n130),
    .overflow(fpu_trans_n131),
    .underflow(fpu_trans_n132),
    .inexact(fpu_trans_n133),
    .invalid(fpu_trans_n134),
    .operation_busy(),
    .operation_done(fpu_trans_n136));
  /* TG68K_FPU.vhd:848:9  */
  tg68k_fpu_converter fpu_converter (
    .clk(clk),
    .nreset(nReset),
    .clkena(clkena),
    .start_conversion(converter_start),
    .source_format(converter_source_format),
    .dest_format(converter_dest_format),
    .data_in(converter_data_in),
    .conversion_done(),
    .conversion_valid(),
    .data_out(),
    .overflow(),
    .underflow(),
    .inexact(),
    .invalid());
  /* TG68K_FPU.vhd:875:9  */
  tg68k_fpu_constantrom fpu_const_rom (
    .clk(clk),
    .nreset(nReset),
    .rom_offset(rom_offset),
    .read_enable(rom_read_enable),
    .constant_out(fpu_const_rom_n173),
    .constant_valid(fpu_const_rom_n174));
  /* TG68K_FPU.vhd:890:9  */
  tg68k_fpu_movem fpu_movem (
    .clk(clk),
    .nreset(nReset),
    .clkena(clkena),
    .start_movem(movem_start),
    .direction(movem_direction),
    .register_mask(movem_register_list),
    .predecrement(movem_predecrement),
    .postincrement(movem_postincrement),
    .fmovem_data_request(fmovem_data_request),
    .fmovem_reg_index(fmovem_reg_index),
    .fmovem_data_write(fmovem_data_write),
    .fmovem_data_in(fmovem_data_in),
    .reg_data_in(movem_reg_data_in),
    .movem_done(movem_done),
    .movem_busy(),
    .fmovem_data_out(\fpu_movem.fmovem_data_out ),
    .reg_address(movem_reg_address),
    .reg_data_out(),
    .reg_write_enable(),
    .address_error(movem_unit_address_error));
  /* TG68K_FPU.vhd:925:9  */
  tg68k_fpu_exception_handler fpu_exception_handler (
    .clk(clk),
    .reset(exception_reset),
    .operation_result(final_result),
    .operation_valid(exception_op_valid),
    .operation_type(exception_op_type),
    .operand_a(alu_operand_a),
    .operand_b(alu_operand_b),
    .overflow_flag(final_overflow),
    .underflow_flag(final_underflow),
    .inexact_flag(final_inexact),
    .invalid_flag(final_invalid),
    .divide_by_zero_flag(alu_divide_by_zero),
    .fpcr(fpcr),
    .fpsr_in(fpsr),
    .fpsr_out(exception_fpsr_out),
    .exception_pending(exception_pending_internal),
    .exception_vector(exception_vector_internal),
    .corrected_result(exception_corrected_result));
  /* TG68K_FPU.vhd:958:28  */
  assign n190 = ~nReset;
  /* TG68K_FPU.vhd:959:48  */
  assign n191 = alu_result_valid | trans_result_valid;
  /* TG68K_FPU.vhd:960:34  */
  assign n193 = {1'b0, alu_operation_code};
  /* TG68K_FPU.vhd:965:102  */
  assign n194 = ~exception_pending_internal;
  /* TG68K_FPU.vhd:965:71  */
  assign n195 = n194 & exception_op_valid;
  /* TG68K_FPU.vhd:965:40  */
  assign n196 = n195 ? exception_fpsr_out : fpsr;
  /* TG68K_FPU.vhd:972:53  */
  assign n197 = exception_pending_internal ? exception_vector_internal : exception_code_internal;
  /* TG68K_FPU.vhd:990:48  */
  assign n202 = fp_registers[639:560]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n204 = n202 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n207 = n204 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:990:48  */
  assign n209 = fp_registers[559:480]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n211 = n209 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n213 = n211 ? 1'b1 : n207;
  /* TG68K_FPU.vhd:990:48  */
  assign n214 = fp_registers[479:400]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n216 = n214 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n218 = n216 ? 1'b1 : n213;
  /* TG68K_FPU.vhd:990:48  */
  assign n219 = fp_registers[399:320]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n221 = n219 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n223 = n221 ? 1'b1 : n218;
  /* TG68K_FPU.vhd:990:48  */
  assign n224 = fp_registers[319:240]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n226 = n224 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n228 = n226 ? 1'b1 : n223;
  /* TG68K_FPU.vhd:990:48  */
  assign n229 = fp_registers[239:160]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n231 = n229 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n233 = n231 ? 1'b1 : n228;
  /* TG68K_FPU.vhd:990:48  */
  assign n234 = fp_registers[159:80]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n236 = n234 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n238 = n236 ? 1'b1 : n233;
  /* TG68K_FPU.vhd:990:48  */
  assign n239 = fp_registers[79:0]; // extract
  /* TG68K_FPU.vhd:990:52  */
  assign n241 = n239 != 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:990:33  */
  assign n243 = n241 ? 1'b1 : n238;
  /* TG68K_FPU.vhd:997:33  */
  assign n245 = fpcr != 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:997:56  */
  assign n247 = fpsr != 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:997:48  */
  assign n248 = n245 | n247;
  /* TG68K_FPU.vhd:997:25  */
  assign n251 = n248 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:1002:73  */
  assign n253 = fpsr[15]; // extract
  /* TG68K_FPU.vhd:1002:66  */
  assign n254 = fpu_exception_i | n253;
  /* TG68K_FPU.vhd:1002:85  */
  assign n255 = fpsr[14]; // extract
  /* TG68K_FPU.vhd:1002:78  */
  assign n256 = n254 | n255;
  /* TG68K_FPU.vhd:1002:97  */
  assign n257 = fpsr[13]; // extract
  /* TG68K_FPU.vhd:1002:90  */
  assign n258 = n256 | n257;
  /* TG68K_FPU.vhd:1002:109  */
  assign n259 = fpsr[12]; // extract
  /* TG68K_FPU.vhd:1002:102  */
  assign n260 = n258 | n259;
  /* TG68K_FPU.vhd:1002:121  */
  assign n261 = fpsr[11]; // extract
  /* TG68K_FPU.vhd:1002:114  */
  assign n262 = n260 | n261;
  /* TG68K_FPU.vhd:1002:133  */
  assign n263 = fpsr[10]; // extract
  /* TG68K_FPU.vhd:1002:126  */
  assign n264 = n262 | n263;
  /* TG68K_FPU.vhd:1002:145  */
  assign n265 = fpsr[9]; // extract
  /* TG68K_FPU.vhd:1002:138  */
  assign n266 = n264 | n265;
  /* TG68K_FPU.vhd:1002:156  */
  assign n267 = fpsr[8]; // extract
  /* TG68K_FPU.vhd:1002:149  */
  assign n268 = n266 | n267;
  /* TG68K_FPU.vhd:1009:56  */
  assign n269 = n268 | fpu_busy_internal;
  /* TG68K_FPU.vhd:1009:96  */
  assign n271 = fpu_state != 4'b0000;
  /* TG68K_FPU.vhd:1009:83  */
  assign n272 = n269 | n271;
  /* TG68K_FPU.vhd:1013:58  */
  assign n273 = n243 | n251;
  /* TG68K_FPU.vhd:1013:25  */
  assign n276 = n273 ? 8'b01100000 : 8'b00000000;
  /* TG68K_FPU.vhd:1013:25  */
  assign n279 = n273 ? 8'b00111100 : 8'b00000100;
  /* TG68K_FPU.vhd:1009:25  */
  assign n281 = n272 ? 8'b11011000 : n276;
  /* TG68K_FPU.vhd:1009:25  */
  assign n283 = n272 ? 8'b11011000 : n279;
  /* TG68K_FPU.vhd:983:17  */
  assign n285 = fpu_just_reset ? 8'b00000000 : n281;
  /* TG68K_FPU.vhd:983:17  */
  assign n287 = fpu_just_reset ? 8'b00000100 : n283;
  /* TG68K_FPU.vhd:1035:27  */
  assign n294 = ~nReset;
  /* TG68K_FPU.vhd:1044:33  */
  assign n297 = fpu_enable ? decoder_operation_code : 7'b0000000;
  /* TG68K_FPU.vhd:1044:33  */
  assign n299 = fpu_enable ? decoder_source_reg : 3'b000;
  /* TG68K_FPU.vhd:1044:33  */
  assign n301 = fpu_enable ? decoder_dest_reg : 3'b000;
  /* TG68K_FPU.vhd:1044:33  */
  assign n303 = fpu_enable ? decoder_source_format : 3'b000;
  /* TG68K_FPU.vhd:1044:33  */
  assign n305 = fpu_enable ? decoder_ea_mode : 3'b000;
  /* TG68K_FPU.vhd:1044:33  */
  assign n307 = fpu_enable ? decoder_ea_register : 3'b000;
  /* TG68K_FPU.vhd:1181:27  */
  assign n743 = ~nReset;
  /* TG68K_FPU.vhd:1234:62  */
  assign n745 = fp_reg_access_valid & fp_reg_write_enable;
  /* TG68K_FPU.vhd:1235:44  */
  assign n746 = {28'b0, fp_reg_write_addr};  //  uext
  /* TG68K_FPU.vhd:1235:84  */
  assign n747 = {1'b0, n746};  //  uext
  /* TG68K_FPU.vhd:1235:84  */
  assign n749 = $signed(n747) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1236:62  */
  assign n752 = 3'b111 - fp_reg_write_addr;
  /* TG68K_FPU.vhd:1234:33  */
  assign n755 = n756 ? n6876 : fp_registers;
  /* TG68K_FPU.vhd:1234:33  */
  assign n756 = n749 & n745;
  /* TG68K_FPU.vhd:1249:76  */
  assign n757 = ~supervisor_mode;
  /* TG68K_FPU.vhd:1263:100  */
  assign n759 = {fsave_frame_format, 24'b000000000000000000000000};
  /* TG68K_FPU.vhd:1249:57  */
  assign n761 = n757 ? 32'b00000000000000000000000000000000 : n759;
  /* TG68K_FPU.vhd:1249:57  */
  assign n763 = n757 ? fpu_done_i : 1'b0;
  /* TG68K_FPU.vhd:1249:57  */
  assign n766 = n757 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:1249:57  */
  assign n769 = n757 ? 4'b1000 : 4'b1001;
  /* TG68K_FPU.vhd:1249:57  */
  assign n771 = n757 ? fsave_frame_format_latched : fsave_frame_format;
  /* TG68K_FPU.vhd:1249:57  */
  assign n773 = n757 ? fsave_counter : 6'b000000;
  /* TG68K_FPU.vhd:1249:57  */
  assign n775 = n757 ? 8'b00100000 : exception_code_internal;
  /* TG68K_FPU.vhd:1268:76  */
  assign n776 = ~supervisor_mode;
  /* TG68K_FPU.vhd:1268:57  */
  assign n778 = n776 ? fpu_done_i : 1'b0;
  /* TG68K_FPU.vhd:1268:57  */
  assign n781 = n776 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:1268:57  */
  assign n784 = n776 ? 4'b1000 : 4'b1010;
  /* TG68K_FPU.vhd:1268:57  */
  assign n786 = n776 ? fsave_counter : 6'b000000;
  /* TG68K_FPU.vhd:1268:57  */
  assign n788 = n776 ? frestore_frame_format : 8'b00000000;
  /* TG68K_FPU.vhd:1268:57  */
  assign n794 = n776 ? 8'b00100000 : exception_code_internal;
  /* TG68K_FPU.vhd:1285:77  */
  assign n795 = command_valid & command_pending;
  /* TG68K_FPU.vhd:1287:65  */
  assign n797 = command_cir == 16'b0000000000000001;
  /* TG68K_FPU.vhd:1289:65  */
  assign n799 = command_cir == 16'b0000000000000010;
  /* TG68K_FPU.vhd:1293:65  */
  assign n801 = command_cir == 16'b0000000000000011;
  assign n802 = {n801, n799, n797};
  /* TG68K_FPU.vhd:1286:57  */
  always @*
    case (n802)
      3'b100: n805 = 1'b1;
      3'b010: n805 = 1'b0;
      3'b001: n805 = fpu_done_i;
      default: n805 = fpu_done_i;
    endcase
  /* TG68K_FPU.vhd:1286:57  */
  always @*
    case (n802)
      3'b100: n808 = 1'b0;
      3'b010: n808 = 1'b0;
      3'b001: n808 = 1'b0;
      default: n808 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:1286:57  */
  always @*
    case (n802)
      3'b100: n812 = 4'b0000;
      3'b010: n812 = 4'b0000;
      3'b001: n812 = 4'b0001;
      default: n812 = fpu_state;
    endcase
  /* TG68K_FPU.vhd:1299:95  */
  assign n813 = ~command_valid;
  /* TG68K_FPU.vhd:1299:77  */
  assign n814 = n813 & command_pending;
  /* TG68K_FPU.vhd:1299:49  */
  assign n817 = n814 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:1299:49  */
  assign n819 = n814 ? 4'b1000 : fpu_state;
  /* TG68K_FPU.vhd:1299:49  */
  assign n821 = n814 ? 8'b00100000 : exception_code_internal;
  /* TG68K_FPU.vhd:1285:49  */
  assign n822 = n795 ? n805 : fpu_done_i;
  /* TG68K_FPU.vhd:1285:49  */
  assign n823 = n795 ? n808 : n817;
  /* TG68K_FPU.vhd:1285:49  */
  assign n824 = n795 ? n812 : n819;
  /* TG68K_FPU.vhd:1285:49  */
  assign n825 = n795 ? exception_code_internal : n821;
  /* TG68K_FPU.vhd:1282:49  */
  assign n826 = fpu_enable ? fpu_done_i : n822;
  /* TG68K_FPU.vhd:1282:49  */
  assign n828 = fpu_enable ? 1'b0 : n823;
  /* TG68K_FPU.vhd:1282:49  */
  assign n830 = fpu_enable ? 4'b0001 : n824;
  /* TG68K_FPU.vhd:1282:49  */
  assign n831 = fpu_enable ? exception_code_internal : n825;
  /* TG68K_FPU.vhd:1266:49  */
  assign n832 = frestore_data_write ? n778 : n826;
  /* TG68K_FPU.vhd:1266:49  */
  assign n833 = frestore_data_write ? n781 : n828;
  /* TG68K_FPU.vhd:1266:49  */
  assign n834 = frestore_data_write ? n784 : n830;
  /* TG68K_FPU.vhd:1266:49  */
  assign n835 = frestore_data_write ? n786 : fsave_counter;
  /* TG68K_FPU.vhd:1266:49  */
  assign n836 = frestore_data_write ? n788 : frestore_frame_format;
  /* TG68K_FPU.vhd:1266:49  */
  assign n839 = frestore_data_write ? n794 : n831;
  /* TG68K_FPU.vhd:1247:49  */
  assign n841 = fsave_data_request ? n761 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1247:49  */
  assign n843 = fsave_data_request ? n763 : n832;
  /* TG68K_FPU.vhd:1247:49  */
  assign n844 = fsave_data_request ? n766 : n833;
  /* TG68K_FPU.vhd:1247:49  */
  assign n846 = fsave_data_request ? n769 : n834;
  /* TG68K_FPU.vhd:1247:49  */
  assign n848 = fsave_data_request ? n771 : fsave_frame_format_latched;
  /* TG68K_FPU.vhd:1247:49  */
  assign n849 = fsave_data_request ? n773 : n835;
  /* TG68K_FPU.vhd:1247:49  */
  assign n850 = fsave_data_request ? frestore_frame_format : n836;
  /* TG68K_FPU.vhd:1247:49  */
  assign n853 = fsave_data_request ? n775 : n839;
  /* TG68K_FPU.vhd:1241:41  */
  assign n855 = fpu_state == 4'b0000;
  /* TG68K_FPU.vhd:1323:65  */
  assign n857 = supervisor_mode ? fpu_exception_i : 1'b1;
  /* TG68K_FPU.vhd:1323:65  */
  assign n859 = supervisor_mode ? restore_privilege_violation : 1'b1;
  /* TG68K_FPU.vhd:1323:65  */
  assign n861 = supervisor_mode ? fpu_state : 4'b1000;
  /* TG68K_FPU.vhd:1323:65  */
  assign n863 = supervisor_mode ? exception_code_internal : 8'b00100000;
  /* TG68K_FPU.vhd:1321:57  */
  assign n865 = decoder_instruction_type == 4'b0110;
  /* TG68K_FPU.vhd:1321:73  */
  assign n867 = decoder_instruction_type == 4'b0111;
  /* TG68K_FPU.vhd:1321:73  */
  assign n868 = n865 | n867;
  /* TG68K_FPU.vhd:1339:133  */
  assign n870 = $unsigned(current_privilege_level) <= $unsigned(3'b001);
  /* TG68K_FPU.vhd:1339:106  */
  assign n871 = supervisor_mode | n870;
  /* TG68K_FPU.vhd:1339:81  */
  assign n873 = n871 ? fpu_exception_i : 1'b1;
  /* TG68K_FPU.vhd:1339:81  */
  assign n875 = n871 ? restore_privilege_violation : 1'b1;
  /* TG68K_FPU.vhd:1339:81  */
  assign n877 = n871 ? fpu_state : 4'b1000;
  /* TG68K_FPU.vhd:1339:81  */
  assign n879 = n871 ? exception_code_internal : 8'b00100000;
  /* TG68K_FPU.vhd:1337:73  */
  assign n881 = extension_word == 16'b1011110000000000;
  /* TG68K_FPU.vhd:1337:86  */
  assign n883 = extension_word == 16'b1001110000000000;
  /* TG68K_FPU.vhd:1337:86  */
  assign n884 = n881 | n883;
  /* TG68K_FPU.vhd:1336:65  */
  always @*
    case (n884)
      1'b1: n885 = n873;
      default: n885 = fpu_exception_i;
    endcase
  /* TG68K_FPU.vhd:1336:65  */
  always @*
    case (n884)
      1'b1: n886 = n875;
      default: n886 = restore_privilege_violation;
    endcase
  /* TG68K_FPU.vhd:1336:65  */
  always @*
    case (n884)
      1'b1: n887 = n877;
      default: n887 = fpu_state;
    endcase
  /* TG68K_FPU.vhd:1336:65  */
  always @*
    case (n884)
      1'b1: n888 = n879;
      default: n888 = exception_code_internal;
    endcase
  /* TG68K_FPU.vhd:1334:57  */
  assign n890 = decoder_instruction_type == 4'b1001;
  /* TG68K_FPU.vhd:1357:92  */
  assign n892 = $unsigned(current_privilege_level) <= $unsigned(3'b001);
  /* TG68K_FPU.vhd:1357:65  */
  assign n894 = n892 ? fpu_exception_i : 1'b1;
  /* TG68K_FPU.vhd:1357:65  */
  assign n896 = n892 ? restore_privilege_violation : 1'b1;
  /* TG68K_FPU.vhd:1357:65  */
  assign n898 = n892 ? fpu_state : 4'b1000;
  /* TG68K_FPU.vhd:1357:65  */
  assign n900 = n892 ? exception_code_internal : 8'b00100000;
  /* TG68K_FPU.vhd:1355:57  */
  assign n902 = decoder_instruction_type == 4'b1000;
  /* TG68K_FPU.vhd:1371:65  */
  assign n904 = fpu_enable ? fpu_exception_i : 1'b1;
  /* TG68K_FPU.vhd:1371:65  */
  assign n906 = fpu_enable ? fpu_state : 4'b1000;
  /* TG68K_FPU.vhd:1371:65  */
  assign n908 = fpu_enable ? exception_code_internal : 8'b00001011;
  assign n909 = {n902, n890, n868};
  /* TG68K_FPU.vhd:1320:49  */
  always @*
    case (n909)
      3'b100: n910 = n894;
      3'b010: n910 = n885;
      3'b001: n910 = n857;
      default: n910 = n904;
    endcase
  /* TG68K_FPU.vhd:1320:49  */
  always @*
    case (n909)
      3'b100: n911 = n896;
      3'b010: n911 = n886;
      3'b001: n911 = n859;
      default: n911 = restore_privilege_violation;
    endcase
  /* TG68K_FPU.vhd:1320:49  */
  always @*
    case (n909)
      3'b100: n912 = n898;
      3'b010: n912 = n887;
      3'b001: n912 = n861;
      default: n912 = n906;
    endcase
  /* TG68K_FPU.vhd:1320:49  */
  always @*
    case (n909)
      3'b100: n913 = n900;
      3'b010: n913 = n888;
      3'b001: n913 = n863;
      default: n913 = n908;
    endcase
  /* TG68K_FPU.vhd:1389:77  */
  assign n915 = decoder_instruction_type != 4'b0101;
  /* TG68K_FPU.vhd:1389:119  */
  assign n917 = decoder_instruction_type != 4'b1001;
  /* TG68K_FPU.vhd:1389:90  */
  assign n918 = n917 & n915;
  /* TG68K_FPU.vhd:1389:49  */
  assign n919 = n918 ? cpu_address_in : fpiar;
  /* TG68K_FPU.vhd:1411:81  */
  assign n920 = ~decoder_valid_instruction;
  /* TG68K_FPU.vhd:1417:72  */
  assign n922 = decoder_instruction_type == 4'b1001;
  /* TG68K_FPU.vhd:480:34  */
  assign n935 = fpsr[31]; // extract
  /* TG68K_FPU.vhd:481:34  */
  assign n937 = fpsr[30]; // extract
  /* TG68K_FPU.vhd:483:34  */
  assign n941 = fpsr[28]; // extract
  /* TG68K_FPU.vhd:486:31  */
  assign n943 = opcode[4:0]; // extract
  /* TG68K_FPU.vhd:487:25  */
  assign n945 = n943 == 5'b00000;
  /* TG68K_FPU.vhd:489:25  */
  assign n947 = n943 == 5'b00001;
  /* TG68K_FPU.vhd:492:55  */
  assign n948 = n941 | n937;
  /* TG68K_FPU.vhd:492:63  */
  assign n949 = n948 | n935;
  /* TG68K_FPU.vhd:492:43  */
  assign n950 = ~n949;
  /* TG68K_FPU.vhd:491:25  */
  assign n952 = n943 == 5'b00010;
  /* TG68K_FPU.vhd:494:64  */
  assign n953 = n941 | n935;
  /* TG68K_FPU.vhd:494:52  */
  assign n954 = ~n953;
  /* TG68K_FPU.vhd:494:48  */
  assign n955 = n937 | n954;
  /* TG68K_FPU.vhd:493:25  */
  assign n957 = n943 == 5'b00011;
  /* TG68K_FPU.vhd:496:65  */
  assign n958 = n941 | n937;
  /* TG68K_FPU.vhd:496:53  */
  assign n959 = ~n958;
  /* TG68K_FPU.vhd:496:48  */
  assign n960 = n935 & n959;
  /* TG68K_FPU.vhd:495:25  */
  assign n962 = n943 == 5'b00100;
  /* TG68K_FPU.vhd:498:62  */
  assign n963 = ~n941;
  /* TG68K_FPU.vhd:498:57  */
  assign n964 = n935 & n963;
  /* TG68K_FPU.vhd:498:48  */
  assign n965 = n937 | n964;
  /* TG68K_FPU.vhd:497:25  */
  assign n967 = n943 == 5'b00101;
  /* TG68K_FPU.vhd:500:44  */
  assign n968 = ~n941;
  /* TG68K_FPU.vhd:500:61  */
  assign n969 = ~n937;
  /* TG68K_FPU.vhd:500:56  */
  assign n970 = n968 & n969;
  /* TG68K_FPU.vhd:499:25  */
  assign n972 = n943 == 5'b00110;
  /* TG68K_FPU.vhd:502:43  */
  assign n973 = ~n941;
  /* TG68K_FPU.vhd:501:25  */
  assign n975 = n943 == 5'b00111;
  /* TG68K_FPU.vhd:503:25  */
  assign n977 = n943 == 5'b01000;
  /* TG68K_FPU.vhd:506:50  */
  assign n978 = n941 | n937;
  /* TG68K_FPU.vhd:505:25  */
  assign n980 = n943 == 5'b01001;
  /* TG68K_FPU.vhd:508:64  */
  assign n981 = n935 | n937;
  /* TG68K_FPU.vhd:508:54  */
  assign n982 = ~n981;
  /* TG68K_FPU.vhd:508:50  */
  assign n983 = n941 | n982;
  /* TG68K_FPU.vhd:507:25  */
  assign n985 = n943 == 5'b01010;
  /* TG68K_FPU.vhd:510:50  */
  assign n986 = n941 | n937;
  /* TG68K_FPU.vhd:510:62  */
  assign n987 = ~n935;
  /* TG68K_FPU.vhd:510:58  */
  assign n988 = n986 | n987;
  /* TG68K_FPU.vhd:509:25  */
  assign n990 = n943 == 5'b01011;
  /* TG68K_FPU.vhd:512:64  */
  assign n991 = ~n937;
  /* TG68K_FPU.vhd:512:59  */
  assign n992 = n935 & n991;
  /* TG68K_FPU.vhd:512:50  */
  assign n993 = n941 | n992;
  /* TG68K_FPU.vhd:511:25  */
  assign n995 = n943 == 5'b01100;
  /* TG68K_FPU.vhd:514:50  */
  assign n996 = n941 | n937;
  /* TG68K_FPU.vhd:514:58  */
  assign n997 = n996 | n935;
  /* TG68K_FPU.vhd:513:25  */
  assign n999 = n943 == 5'b01101;
  /* TG68K_FPU.vhd:516:43  */
  assign n1000 = ~n937;
  /* TG68K_FPU.vhd:515:25  */
  assign n1002 = n943 == 5'b01110;
  /* TG68K_FPU.vhd:517:25  */
  assign n1004 = n943 == 5'b01111;
  assign n1005 = {n1004, n1002, n999, n995, n990, n985, n980, n977, n975, n972, n967, n962, n957, n952, n947, n945};
  /* TG68K_FPU.vhd:486:17  */
  always @*
    case (n1005)
      16'b1000000000000000: n1009 = 1'b1;
      16'b0100000000000000: n1009 = n1000;
      16'b0010000000000000: n1009 = n997;
      16'b0001000000000000: n1009 = n993;
      16'b0000100000000000: n1009 = n988;
      16'b0000010000000000: n1009 = n983;
      16'b0000001000000000: n1009 = n978;
      16'b0000000100000000: n1009 = n941;
      16'b0000000010000000: n1009 = n973;
      16'b0000000001000000: n1009 = n970;
      16'b0000000000100000: n1009 = n965;
      16'b0000000000010000: n1009 = n960;
      16'b0000000000001000: n1009 = n955;
      16'b0000000000000100: n1009 = n950;
      16'b0000000000000010: n1009 = n937;
      16'b0000000000000001: n1009 = 1'b0;
      default: n1009 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:1425:110  */
  assign n1012 = cpu_data_in - 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:1420:49  */
  assign n1014 = n1009 ? 32'b00000000000000000000000000000001 : n1012;
  /* TG68K_FPU.vhd:1431:72  */
  assign n1016 = decoder_instruction_type == 4'b0101;
  /* TG68K_FPU.vhd:480:34  */
  assign n1029 = fpsr[31]; // extract
  /* TG68K_FPU.vhd:481:34  */
  assign n1031 = fpsr[30]; // extract
  /* TG68K_FPU.vhd:483:34  */
  assign n1035 = fpsr[28]; // extract
  /* TG68K_FPU.vhd:486:31  */
  assign n1037 = opcode[4:0]; // extract
  /* TG68K_FPU.vhd:487:25  */
  assign n1039 = n1037 == 5'b00000;
  /* TG68K_FPU.vhd:489:25  */
  assign n1041 = n1037 == 5'b00001;
  /* TG68K_FPU.vhd:492:55  */
  assign n1042 = n1035 | n1031;
  /* TG68K_FPU.vhd:492:63  */
  assign n1043 = n1042 | n1029;
  /* TG68K_FPU.vhd:492:43  */
  assign n1044 = ~n1043;
  /* TG68K_FPU.vhd:491:25  */
  assign n1046 = n1037 == 5'b00010;
  /* TG68K_FPU.vhd:494:64  */
  assign n1047 = n1035 | n1029;
  /* TG68K_FPU.vhd:494:52  */
  assign n1048 = ~n1047;
  /* TG68K_FPU.vhd:494:48  */
  assign n1049 = n1031 | n1048;
  /* TG68K_FPU.vhd:493:25  */
  assign n1051 = n1037 == 5'b00011;
  /* TG68K_FPU.vhd:496:65  */
  assign n1052 = n1035 | n1031;
  /* TG68K_FPU.vhd:496:53  */
  assign n1053 = ~n1052;
  /* TG68K_FPU.vhd:496:48  */
  assign n1054 = n1029 & n1053;
  /* TG68K_FPU.vhd:495:25  */
  assign n1056 = n1037 == 5'b00100;
  /* TG68K_FPU.vhd:498:62  */
  assign n1057 = ~n1035;
  /* TG68K_FPU.vhd:498:57  */
  assign n1058 = n1029 & n1057;
  /* TG68K_FPU.vhd:498:48  */
  assign n1059 = n1031 | n1058;
  /* TG68K_FPU.vhd:497:25  */
  assign n1061 = n1037 == 5'b00101;
  /* TG68K_FPU.vhd:500:44  */
  assign n1062 = ~n1035;
  /* TG68K_FPU.vhd:500:61  */
  assign n1063 = ~n1031;
  /* TG68K_FPU.vhd:500:56  */
  assign n1064 = n1062 & n1063;
  /* TG68K_FPU.vhd:499:25  */
  assign n1066 = n1037 == 5'b00110;
  /* TG68K_FPU.vhd:502:43  */
  assign n1067 = ~n1035;
  /* TG68K_FPU.vhd:501:25  */
  assign n1069 = n1037 == 5'b00111;
  /* TG68K_FPU.vhd:503:25  */
  assign n1071 = n1037 == 5'b01000;
  /* TG68K_FPU.vhd:506:50  */
  assign n1072 = n1035 | n1031;
  /* TG68K_FPU.vhd:505:25  */
  assign n1074 = n1037 == 5'b01001;
  /* TG68K_FPU.vhd:508:64  */
  assign n1075 = n1029 | n1031;
  /* TG68K_FPU.vhd:508:54  */
  assign n1076 = ~n1075;
  /* TG68K_FPU.vhd:508:50  */
  assign n1077 = n1035 | n1076;
  /* TG68K_FPU.vhd:507:25  */
  assign n1079 = n1037 == 5'b01010;
  /* TG68K_FPU.vhd:510:50  */
  assign n1080 = n1035 | n1031;
  /* TG68K_FPU.vhd:510:62  */
  assign n1081 = ~n1029;
  /* TG68K_FPU.vhd:510:58  */
  assign n1082 = n1080 | n1081;
  /* TG68K_FPU.vhd:509:25  */
  assign n1084 = n1037 == 5'b01011;
  /* TG68K_FPU.vhd:512:64  */
  assign n1085 = ~n1031;
  /* TG68K_FPU.vhd:512:59  */
  assign n1086 = n1029 & n1085;
  /* TG68K_FPU.vhd:512:50  */
  assign n1087 = n1035 | n1086;
  /* TG68K_FPU.vhd:511:25  */
  assign n1089 = n1037 == 5'b01100;
  /* TG68K_FPU.vhd:514:50  */
  assign n1090 = n1035 | n1031;
  /* TG68K_FPU.vhd:514:58  */
  assign n1091 = n1090 | n1029;
  /* TG68K_FPU.vhd:513:25  */
  assign n1093 = n1037 == 5'b01101;
  /* TG68K_FPU.vhd:516:43  */
  assign n1094 = ~n1031;
  /* TG68K_FPU.vhd:515:25  */
  assign n1096 = n1037 == 5'b01110;
  /* TG68K_FPU.vhd:517:25  */
  assign n1098 = n1037 == 5'b01111;
  assign n1099 = {n1098, n1096, n1093, n1089, n1084, n1079, n1074, n1071, n1069, n1066, n1061, n1056, n1051, n1046, n1041, n1039};
  /* TG68K_FPU.vhd:486:17  */
  always @*
    case (n1099)
      16'b1000000000000000: n1103 = 1'b1;
      16'b0100000000000000: n1103 = n1094;
      16'b0010000000000000: n1103 = n1091;
      16'b0001000000000000: n1103 = n1087;
      16'b0000100000000000: n1103 = n1082;
      16'b0000010000000000: n1103 = n1077;
      16'b0000001000000000: n1103 = n1072;
      16'b0000000100000000: n1103 = n1035;
      16'b0000000010000000: n1103 = n1067;
      16'b0000000001000000: n1103 = n1064;
      16'b0000000000100000: n1103 = n1059;
      16'b0000000000010000: n1103 = n1054;
      16'b0000000000001000: n1103 = n1049;
      16'b0000000000000100: n1103 = n1044;
      16'b0000000000000010: n1103 = n1031;
      16'b0000000000000001: n1103 = 1'b0;
      default: n1103 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:1434:49  */
  assign n1107 = n1103 ? 32'b00000000000000000000000000000001 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1442:72  */
  assign n1109 = decoder_instruction_type == 4'b1000;
  /* TG68K_FPU.vhd:480:34  */
  assign n1122 = fpsr[31]; // extract
  /* TG68K_FPU.vhd:481:34  */
  assign n1124 = fpsr[30]; // extract
  /* TG68K_FPU.vhd:483:34  */
  assign n1128 = fpsr[28]; // extract
  /* TG68K_FPU.vhd:486:31  */
  assign n1130 = opcode[4:0]; // extract
  /* TG68K_FPU.vhd:487:25  */
  assign n1132 = n1130 == 5'b00000;
  /* TG68K_FPU.vhd:489:25  */
  assign n1134 = n1130 == 5'b00001;
  /* TG68K_FPU.vhd:492:55  */
  assign n1135 = n1128 | n1124;
  /* TG68K_FPU.vhd:492:63  */
  assign n1136 = n1135 | n1122;
  /* TG68K_FPU.vhd:492:43  */
  assign n1137 = ~n1136;
  /* TG68K_FPU.vhd:491:25  */
  assign n1139 = n1130 == 5'b00010;
  /* TG68K_FPU.vhd:494:64  */
  assign n1140 = n1128 | n1122;
  /* TG68K_FPU.vhd:494:52  */
  assign n1141 = ~n1140;
  /* TG68K_FPU.vhd:494:48  */
  assign n1142 = n1124 | n1141;
  /* TG68K_FPU.vhd:493:25  */
  assign n1144 = n1130 == 5'b00011;
  /* TG68K_FPU.vhd:496:65  */
  assign n1145 = n1128 | n1124;
  /* TG68K_FPU.vhd:496:53  */
  assign n1146 = ~n1145;
  /* TG68K_FPU.vhd:496:48  */
  assign n1147 = n1122 & n1146;
  /* TG68K_FPU.vhd:495:25  */
  assign n1149 = n1130 == 5'b00100;
  /* TG68K_FPU.vhd:498:62  */
  assign n1150 = ~n1128;
  /* TG68K_FPU.vhd:498:57  */
  assign n1151 = n1122 & n1150;
  /* TG68K_FPU.vhd:498:48  */
  assign n1152 = n1124 | n1151;
  /* TG68K_FPU.vhd:497:25  */
  assign n1154 = n1130 == 5'b00101;
  /* TG68K_FPU.vhd:500:44  */
  assign n1155 = ~n1128;
  /* TG68K_FPU.vhd:500:61  */
  assign n1156 = ~n1124;
  /* TG68K_FPU.vhd:500:56  */
  assign n1157 = n1155 & n1156;
  /* TG68K_FPU.vhd:499:25  */
  assign n1159 = n1130 == 5'b00110;
  /* TG68K_FPU.vhd:502:43  */
  assign n1160 = ~n1128;
  /* TG68K_FPU.vhd:501:25  */
  assign n1162 = n1130 == 5'b00111;
  /* TG68K_FPU.vhd:503:25  */
  assign n1164 = n1130 == 5'b01000;
  /* TG68K_FPU.vhd:506:50  */
  assign n1165 = n1128 | n1124;
  /* TG68K_FPU.vhd:505:25  */
  assign n1167 = n1130 == 5'b01001;
  /* TG68K_FPU.vhd:508:64  */
  assign n1168 = n1122 | n1124;
  /* TG68K_FPU.vhd:508:54  */
  assign n1169 = ~n1168;
  /* TG68K_FPU.vhd:508:50  */
  assign n1170 = n1128 | n1169;
  /* TG68K_FPU.vhd:507:25  */
  assign n1172 = n1130 == 5'b01010;
  /* TG68K_FPU.vhd:510:50  */
  assign n1173 = n1128 | n1124;
  /* TG68K_FPU.vhd:510:62  */
  assign n1174 = ~n1122;
  /* TG68K_FPU.vhd:510:58  */
  assign n1175 = n1173 | n1174;
  /* TG68K_FPU.vhd:509:25  */
  assign n1177 = n1130 == 5'b01011;
  /* TG68K_FPU.vhd:512:64  */
  assign n1178 = ~n1124;
  /* TG68K_FPU.vhd:512:59  */
  assign n1179 = n1122 & n1178;
  /* TG68K_FPU.vhd:512:50  */
  assign n1180 = n1128 | n1179;
  /* TG68K_FPU.vhd:511:25  */
  assign n1182 = n1130 == 5'b01100;
  /* TG68K_FPU.vhd:514:50  */
  assign n1183 = n1128 | n1124;
  /* TG68K_FPU.vhd:514:58  */
  assign n1184 = n1183 | n1122;
  /* TG68K_FPU.vhd:513:25  */
  assign n1186 = n1130 == 5'b01101;
  /* TG68K_FPU.vhd:516:43  */
  assign n1187 = ~n1124;
  /* TG68K_FPU.vhd:515:25  */
  assign n1189 = n1130 == 5'b01110;
  /* TG68K_FPU.vhd:517:25  */
  assign n1191 = n1130 == 5'b01111;
  assign n1192 = {n1191, n1189, n1186, n1182, n1177, n1172, n1167, n1164, n1162, n1159, n1154, n1149, n1144, n1139, n1134, n1132};
  /* TG68K_FPU.vhd:486:17  */
  always @*
    case (n1192)
      16'b1000000000000000: n1196 = 1'b1;
      16'b0100000000000000: n1196 = n1187;
      16'b0010000000000000: n1196 = n1184;
      16'b0001000000000000: n1196 = n1180;
      16'b0000100000000000: n1196 = n1175;
      16'b0000010000000000: n1196 = n1170;
      16'b0000001000000000: n1196 = n1165;
      16'b0000000100000000: n1196 = n1128;
      16'b0000000010000000: n1196 = n1160;
      16'b0000000001000000: n1196 = n1157;
      16'b0000000000100000: n1196 = n1152;
      16'b0000000000010000: n1196 = n1147;
      16'b0000000000001000: n1196 = n1142;
      16'b0000000000000100: n1196 = n1137;
      16'b0000000000000010: n1196 = n1124;
      16'b0000000000000001: n1196 = 1'b0;
      default: n1196 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:1445:49  */
  assign n1200 = n1196 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:1445:49  */
  assign n1202 = n1196 ? 1'b1 : n910;
  /* TG68K_FPU.vhd:1445:49  */
  assign n1205 = n1196 ? 4'b1000 : 4'b0000;
  /* TG68K_FPU.vhd:1445:49  */
  assign n1207 = n1196 ? 8'b00000111 : n913;
  /* TG68K_FPU.vhd:1457:72  */
  assign n1209 = decoder_instruction_type == 4'b0000;
  /* TG68K_FPU.vhd:1458:74  */
  assign n1211 = decoder_operation_code == 7'b0111010;
  /* TG68K_FPU.vhd:1457:87  */
  assign n1212 = n1211 & n1209;
  /* TG68K_FPU.vhd:1459:67  */
  assign n1214 = decoder_ea_mode == 3'b000;
  /* TG68K_FPU.vhd:1458:84  */
  assign n1215 = n1214 & n1212;
  /* TG68K_FPU.vhd:1467:79  */
  assign n1216 = cpu_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:1467:92  */
  assign n1218 = n1216 == 8'b00000000;
  /* TG68K_FPU.vhd:1469:82  */
  assign n1220 = cpu_data_in[7]; // extract
  /* TG68K_FPU.vhd:1469:65  */
  assign n1223 = n1220 ? 4'b1000 : 4'b0000;
  /* TG68K_FPU.vhd:1467:65  */
  assign n1224 = n1218 ? 4'b0100 : n1223;
  /* TG68K_FPU.vhd:1464:57  */
  assign n1226 = decoder_source_format == 3'b110;
  /* TG68K_FPU.vhd:1476:79  */
  assign n1227 = cpu_data_in[15:0]; // extract
  /* TG68K_FPU.vhd:1476:93  */
  assign n1229 = n1227 == 16'b0000000000000000;
  /* TG68K_FPU.vhd:1478:82  */
  assign n1231 = cpu_data_in[15]; // extract
  /* TG68K_FPU.vhd:1478:65  */
  assign n1234 = n1231 ? 4'b1000 : 4'b0000;
  /* TG68K_FPU.vhd:1476:65  */
  assign n1235 = n1229 ? 4'b0100 : n1234;
  /* TG68K_FPU.vhd:1474:57  */
  assign n1237 = decoder_source_format == 3'b100;
  /* TG68K_FPU.vhd:1485:80  */
  assign n1239 = cpu_data_in == 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1487:82  */
  assign n1241 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:1487:65  */
  assign n1244 = n1241 ? 4'b1000 : 4'b0000;
  /* TG68K_FPU.vhd:1485:65  */
  assign n1245 = n1239 ? 4'b0100 : n1244;
  /* TG68K_FPU.vhd:1483:57  */
  assign n1247 = decoder_source_format == 3'b000;
  assign n1249 = {n1247, n1237, n1226};
  /* TG68K_FPU.vhd:1463:49  */
  always @*
    case (n1249)
      3'b100: n1250 = n1245;
      3'b010: n1250 = n1235;
      3'b001: n1250 = n1224;
      default: n1250 = 4'b0001;
    endcase
  /* TG68K_FPU.vhd:1499:72  */
  assign n1252 = decoder_instruction_type == 4'b0000;
  /* TG68K_FPU.vhd:1500:75  */
  assign n1254 = decoder_operation_code == 7'b0011000;
  /* TG68K_FPU.vhd:1500:111  */
  assign n1256 = decoder_operation_code == 7'b0011010;
  /* TG68K_FPU.vhd:1500:85  */
  assign n1257 = n1254 | n1256;
  /* TG68K_FPU.vhd:1500:147  */
  assign n1259 = decoder_operation_code == 7'b0000000;
  /* TG68K_FPU.vhd:1500:121  */
  assign n1260 = n1257 | n1259;
  /* TG68K_FPU.vhd:1500:184  */
  assign n1262 = decoder_operation_code == 7'b1000001;
  /* TG68K_FPU.vhd:1500:158  */
  assign n1263 = n1260 | n1262;
  /* TG68K_FPU.vhd:1499:87  */
  assign n1264 = n1263 & n1252;
  /* TG68K_FPU.vhd:1501:70  */
  assign n1266 = decoder_source_reg != 3'b111;
  /* TG68K_FPU.vhd:1500:198  */
  assign n1267 = n1266 & n1264;
  /* TG68K_FPU.vhd:1507:68  */
  assign n1268 = {28'b0, decoder_source_reg};  //  uext
  /* TG68K_FPU.vhd:1507:109  */
  assign n1269 = {1'b0, n1268};  //  uext
  /* TG68K_FPU.vhd:1507:109  */
  assign n1271 = $signed(n1269) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1507:118  */
  assign n1272 = {28'b0, decoder_dest_reg};  //  uext
  /* TG68K_FPU.vhd:1507:157  */
  assign n1273 = {1'b0, n1272};  //  uext
  /* TG68K_FPU.vhd:1507:157  */
  assign n1275 = $signed(n1273) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1507:114  */
  assign n1276 = n1275 & n1271;
  /* TG68K_FPU.vhd:1510:113  */
  assign n1279 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1510:154  */
  assign n1281 = fp_registers[n6879 + 0 +: 79]; //(dyn_extract)
  /* TG68K_FPU.vhd:1510:98  */
  assign n1283 = {1'b0, n1281};
  /* TG68K_FPU.vhd:1507:65  */
  assign n1285 = n1276 ? n910 : 1'b1;
  /* TG68K_FPU.vhd:1507:65  */
  assign n1287 = n1276 ? 1'b1 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:1507:65  */
  assign n1288 = n1276 ? decoder_dest_reg : fp_reg_write_addr;
  /* TG68K_FPU.vhd:1507:65  */
  assign n1289 = n1276 ? n1283 : fp_reg_write_data;
  /* TG68K_FPU.vhd:1507:65  */
  assign n1292 = n1276 ? 1'b1 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:1507:65  */
  assign n1294 = n1276 ? n912 : 4'b1000;
  /* TG68K_FPU.vhd:1507:65  */
  assign n1296 = n1276 ? n913 : 8'b00010100;
  /* TG68K_FPU.vhd:1504:57  */
  assign n1298 = decoder_operation_code == 7'b0011000;
  /* TG68K_FPU.vhd:1522:68  */
  assign n1299 = {28'b0, decoder_source_reg};  //  uext
  /* TG68K_FPU.vhd:1522:109  */
  assign n1300 = {1'b0, n1299};  //  uext
  /* TG68K_FPU.vhd:1522:109  */
  assign n1302 = $signed(n1300) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1522:118  */
  assign n1303 = {28'b0, decoder_dest_reg};  //  uext
  /* TG68K_FPU.vhd:1522:157  */
  assign n1304 = {1'b0, n1303};  //  uext
  /* TG68K_FPU.vhd:1522:157  */
  assign n1306 = $signed(n1304) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1522:114  */
  assign n1307 = n1306 & n1302;
  /* TG68K_FPU.vhd:1525:111  */
  assign n1310 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1525:94  */
  assign n1313 = ~n6884;
  /* TG68K_FPU.vhd:1526:126  */
  assign n1316 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1526:167  */
  assign n1318 = fp_registers[n6887 + 0 +: 79]; //(dyn_extract)
  /* TG68K_FPU.vhd:1525:157  */
  assign n1319 = {n1313, n1318};
  /* TG68K_FPU.vhd:1522:65  */
  assign n1321 = n1307 ? n910 : 1'b1;
  /* TG68K_FPU.vhd:1522:65  */
  assign n1323 = n1307 ? 1'b1 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:1522:65  */
  assign n1324 = n1307 ? decoder_dest_reg : fp_reg_write_addr;
  /* TG68K_FPU.vhd:1522:65  */
  assign n1325 = n1307 ? n1319 : fp_reg_write_data;
  /* TG68K_FPU.vhd:1522:65  */
  assign n1328 = n1307 ? 1'b1 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:1522:65  */
  assign n1330 = n1307 ? n912 : 4'b1000;
  /* TG68K_FPU.vhd:1522:65  */
  assign n1332 = n1307 ? n913 : 8'b00010100;
  /* TG68K_FPU.vhd:1519:57  */
  assign n1334 = decoder_operation_code == 7'b0011010;
  /* TG68K_FPU.vhd:1538:68  */
  assign n1335 = {28'b0, decoder_source_reg};  //  uext
  /* TG68K_FPU.vhd:1538:109  */
  assign n1336 = {1'b0, n1335};  //  uext
  /* TG68K_FPU.vhd:1538:109  */
  assign n1338 = $signed(n1336) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1538:118  */
  assign n1339 = {28'b0, decoder_dest_reg};  //  uext
  /* TG68K_FPU.vhd:1538:157  */
  assign n1340 = {1'b0, n1339};  //  uext
  /* TG68K_FPU.vhd:1538:157  */
  assign n1342 = $signed(n1340) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1538:114  */
  assign n1343 = n1342 & n1338;
  /* TG68K_FPU.vhd:1541:107  */
  assign n1346 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1538:65  */
  assign n1350 = n1343 ? n910 : 1'b1;
  /* TG68K_FPU.vhd:1538:65  */
  assign n1352 = n1343 ? 1'b1 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:1538:65  */
  assign n1353 = n1343 ? decoder_dest_reg : fp_reg_write_addr;
  /* TG68K_FPU.vhd:1538:65  */
  assign n1354 = n1343 ? n6888 : fp_reg_write_data;
  /* TG68K_FPU.vhd:1538:65  */
  assign n1357 = n1343 ? 1'b1 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:1538:65  */
  assign n1359 = n1343 ? n912 : 4'b1000;
  /* TG68K_FPU.vhd:1538:65  */
  assign n1361 = n1343 ? n913 : 8'b00010100;
  /* TG68K_FPU.vhd:1535:57  */
  assign n1363 = decoder_operation_code == 7'b0000000;
  /* TG68K_FPU.vhd:1552:98  */
  assign n1365 = {decoder_source_reg, 4'b0000};
  /* TG68K_FPU.vhd:1550:57  */
  assign n1367 = decoder_operation_code == 7'b1000001;
  /* TG68K_FPU.vhd:1560:76  */
  assign n1368 = opcode[5:0]; // extract
  /* TG68K_FPU.vhd:1560:89  */
  assign n1370 = n1368 == 6'b000001;
  /* TG68K_FPU.vhd:1560:108  */
  assign n1371 = fpsr[29]; // extract
  /* TG68K_FPU.vhd:1560:100  */
  assign n1372 = n1371 & n1370;
  /* TG68K_FPU.vhd:1561:76  */
  assign n1373 = opcode[5:0]; // extract
  /* TG68K_FPU.vhd:1561:89  */
  assign n1375 = n1373 == 6'b001110;
  /* TG68K_FPU.vhd:1561:108  */
  assign n1376 = fpsr[29]; // extract
  /* TG68K_FPU.vhd:1561:113  */
  assign n1377 = ~n1376;
  /* TG68K_FPU.vhd:1561:100  */
  assign n1378 = n1377 & n1375;
  /* TG68K_FPU.vhd:1560:120  */
  assign n1379 = n1372 | n1378;
  /* TG68K_FPU.vhd:1562:76  */
  assign n1380 = opcode[5:0]; // extract
  /* TG68K_FPU.vhd:1562:89  */
  assign n1382 = n1380 == 6'b010010;
  /* TG68K_FPU.vhd:1562:108  */
  assign n1383 = fpsr[28]; // extract
  /* TG68K_FPU.vhd:1562:100  */
  assign n1384 = n1383 & n1382;
  /* TG68K_FPU.vhd:1561:120  */
  assign n1385 = n1379 | n1384;
  /* TG68K_FPU.vhd:1563:76  */
  assign n1386 = opcode[5:0]; // extract
  /* TG68K_FPU.vhd:1563:89  */
  assign n1388 = n1386 == 6'b010011;
  /* TG68K_FPU.vhd:1563:108  */
  assign n1389 = fpsr[29]; // extract
  /* TG68K_FPU.vhd:1563:100  */
  assign n1390 = n1389 & n1388;
  /* TG68K_FPU.vhd:1562:120  */
  assign n1391 = n1385 | n1390;
  /* TG68K_FPU.vhd:1564:76  */
  assign n1392 = opcode[5:0]; // extract
  /* TG68K_FPU.vhd:1564:89  */
  assign n1394 = n1392 == 6'b010100;
  /* TG68K_FPU.vhd:1564:108  */
  assign n1395 = fpsr[30]; // extract
  /* TG68K_FPU.vhd:1564:100  */
  assign n1396 = n1395 & n1394;
  /* TG68K_FPU.vhd:1563:120  */
  assign n1397 = n1391 | n1396;
  /* TG68K_FPU.vhd:1565:76  */
  assign n1398 = opcode[5:0]; // extract
  /* TG68K_FPU.vhd:1565:89  */
  assign n1400 = n1398 == 6'b010101;
  /* TG68K_FPU.vhd:1565:109  */
  assign n1401 = fpsr[30]; // extract
  /* TG68K_FPU.vhd:1565:127  */
  assign n1402 = fpsr[29]; // extract
  /* TG68K_FPU.vhd:1565:120  */
  assign n1403 = n1401 | n1402;
  /* TG68K_FPU.vhd:1565:100  */
  assign n1404 = n1403 & n1400;
  /* TG68K_FPU.vhd:1564:120  */
  assign n1405 = n1397 | n1404;
  /* TG68K_FPU.vhd:1560:65  */
  assign n1408 = n1405 ? 32'b00000000000000000000000011111111 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1557:57  */
  assign n1410 = decoder_operation_code == 7'b1000010;
  assign n1411 = {n1410, n1367, n1363, n1334, n1298};
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1413 = n1408;
      5'b01000: n1413 = 32'b00000000000000000000000000000000;
      5'b00100: n1413 = 32'b00000000000000000000000000000000;
      5'b00010: n1413 = 32'b00000000000000000000000000000000;
      5'b00001: n1413 = 32'b00000000000000000000000000000000;
      default: n1413 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1416 = 1'b1;
      5'b01000: n1416 = 1'b0;
      5'b00100: n1416 = 1'b0;
      5'b00010: n1416 = 1'b0;
      5'b00001: n1416 = 1'b0;
      default: n1416 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1417 = n910;
      5'b01000: n1417 = n910;
      5'b00100: n1417 = n1350;
      5'b00010: n1417 = n1321;
      5'b00001: n1417 = n1285;
      default: n1417 = n910;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1418 = fp_reg_write_enable;
      5'b01000: n1418 = fp_reg_write_enable;
      5'b00100: n1418 = n1352;
      5'b00010: n1418 = n1323;
      5'b00001: n1418 = n1287;
      default: n1418 = fp_reg_write_enable;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1419 = fp_reg_write_addr;
      5'b01000: n1419 = fp_reg_write_addr;
      5'b00100: n1419 = n1353;
      5'b00010: n1419 = n1324;
      5'b00001: n1419 = n1288;
      default: n1419 = fp_reg_write_addr;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1420 = fp_reg_write_data;
      5'b01000: n1420 = fp_reg_write_data;
      5'b00100: n1420 = n1354;
      5'b00010: n1420 = n1325;
      5'b00001: n1420 = n1289;
      default: n1420 = fp_reg_write_data;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1422 = fp_reg_access_valid;
      5'b01000: n1422 = fp_reg_access_valid;
      5'b00100: n1422 = n1357;
      5'b00010: n1422 = n1328;
      5'b00001: n1422 = n1292;
      default: n1422 = fp_reg_access_valid;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1425 = 4'b0000;
      5'b01000: n1425 = 4'b0110;
      5'b00100: n1425 = n1359;
      5'b00010: n1425 = n1330;
      5'b00001: n1425 = n1294;
      default: n1425 = n912;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1426 = n913;
      5'b01000: n1426 = n913;
      5'b00100: n1426 = n1361;
      5'b00010: n1426 = n1332;
      5'b00001: n1426 = n1296;
      default: n1426 = n913;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1427 = rom_offset;
      5'b01000: n1427 = n1365;
      5'b00100: n1427 = rom_offset;
      5'b00010: n1427 = rom_offset;
      5'b00001: n1427 = rom_offset;
      default: n1427 = rom_offset;
    endcase
  /* TG68K_FPU.vhd:1503:49  */
  always @*
    case (n1411)
      5'b10000: n1429 = rom_read_enable;
      5'b01000: n1429 = 1'b1;
      5'b00100: n1429 = rom_read_enable;
      5'b00010: n1429 = rom_read_enable;
      5'b00001: n1429 = rom_read_enable;
      default: n1429 = rom_read_enable;
    endcase
  /* TG68K_FPU.vhd:1576:75  */
  assign n1431 = decoder_operation_code != 7'b1000001;
  /* TG68K_FPU.vhd:1576:116  */
  assign n1433 = decoder_operation_code != 7'b1000010;
  /* TG68K_FPU.vhd:1576:89  */
  assign n1434 = n1433 & n1431;
  /* TG68K_FPU.vhd:1578:101  */
  assign n1438 = 3'b111 - decoder_dest_reg;
  /* TG68K_FPU.vhd:550:33  */
  assign n1446 = n6889[79]; // extract
  /* TG68K_FPU.vhd:551:37  */
  assign n1448 = n6889[78:64]; // extract
  /* TG68K_FPU.vhd:552:37  */
  assign n1450 = n6889[63:0]; // extract
  /* TG68K_FPU.vhd:558:29  */
  assign n1454 = n1448 == 15'b111111111111111;
  /* TG68K_FPU.vhd:560:36  */
  assign n1455 = n6889[63]; // extract
  /* TG68K_FPU.vhd:560:41  */
  assign n1456 = ~n1455;
  /* TG68K_FPU.vhd:560:58  */
  assign n1457 = n6889[62:0]; // extract
  /* TG68K_FPU.vhd:560:72  */
  assign n1459 = n1457 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:560:47  */
  assign n1460 = n1456 | n1459;
  assign n1463 = n1452[0]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n1464 = n1460 ? 1'b1 : n1463;
  assign n1465 = n1452[1]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n1466 = n1460 ? n1465 : 1'b1;
  assign n1467 = n1452[3]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n1468 = n1460 ? n1467 : n1446;
  /* TG68K_FPU.vhd:568:32  */
  assign n1470 = n1448 == 15'b000000000000000;
  /* TG68K_FPU.vhd:568:68  */
  assign n1472 = n1450 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:568:55  */
  assign n1473 = n1472 & n1470;
  assign n1475 = {n1446, 1'b1};
  assign n1476 = n1475[0]; // extract
  assign n1477 = n1452[2]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n1478 = n1473 ? n1476 : n1477;
  assign n1479 = n1475[1]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n1480 = n1473 ? n1479 : n1446;
  assign n1481 = {n1480, n1478};
  assign n1482 = {n1466, n1464};
  assign n1483 = n1452[1:0]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n1484 = n1454 ? n1482 : n1483;
  assign n1485 = n1481[0]; // extract
  assign n1486 = n1452[2]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n1487 = n1454 ? n1486 : n1485;
  assign n1488 = n1481[1]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n1489 = n1454 ? n1468 : n1488;
  /* TG68K_FPU.vhd:1576:49  */
  assign n1493 = n1434 ? 1'b1 : n1416;
  assign n1494 = {n1489, n1487, n1484};
  assign n1495 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:1576:49  */
  assign n1496 = n1434 ? n1494 : n1495;
  /* TG68K_FPU.vhd:1576:49  */
  assign n1498 = n1434 ? 4'b0000 : n1425;
  /* TG68K_FPU.vhd:1582:72  */
  assign n1500 = decoder_instruction_type == 4'b0011;
  /* TG68K_FPU.vhd:1585:59  */
  assign n1501 = opcode[15:8]; // extract
  /* TG68K_FPU.vhd:1585:73  */
  assign n1503 = n1501 != 8'b11110010;
  /* TG68K_FPU.vhd:1586:67  */
  assign n1504 = extension_word[15:14]; // extract
  /* TG68K_FPU.vhd:1586:82  */
  assign n1506 = n1504 != 2'b11;
  /* TG68K_FPU.vhd:1585:83  */
  assign n1507 = n1503 | n1506;
  /* TG68K_FPU.vhd:1587:67  */
  assign n1508 = extension_word[12:8]; // extract
  /* TG68K_FPU.vhd:1587:81  */
  assign n1510 = n1508 != 5'b00000;
  /* TG68K_FPU.vhd:1586:91  */
  assign n1511 = n1507 | n1510;
  /* TG68K_FPU.vhd:1588:67  */
  assign n1512 = extension_word[7:0]; // extract
  /* TG68K_FPU.vhd:1588:80  */
  assign n1514 = n1512 == 8'b00000000;
  /* TG68K_FPU.vhd:1587:93  */
  assign n1515 = n1511 | n1514;
  /* TG68K_FPU.vhd:1595:94  */
  assign n1516 = extension_word[7:0]; // extract
  /* TG68K_FPU.vhd:1596:90  */
  assign n1517 = extension_word[13]; // extract
  /* TG68K_FPU.vhd:1599:57  */
  assign n1519 = ea_mode == 3'b010;
  /* TG68K_FPU.vhd:1602:57  */
  assign n1521 = ea_mode == 3'b011;
  /* TG68K_FPU.vhd:1606:57  */
  assign n1523 = ea_mode == 3'b100;
  /* TG68K_FPU.vhd:1610:57  */
  assign n1525 = ea_mode == 3'b101;
  /* TG68K_FPU.vhd:1614:57  */
  assign n1532 = ea_mode == 3'b110;
  /* TG68K_FPU.vhd:1625:73  */
  assign n1534 = ea_register == 3'b000;
  /* TG68K_FPU.vhd:1629:73  */
  assign n1536 = ea_register == 3'b001;
  /* TG68K_FPU.vhd:1633:73  */
  assign n1538 = ea_register == 3'b010;
  /* TG68K_FPU.vhd:1636:73  */
  assign n1540 = ea_register == 3'b011;
  /* TG68K_FPU.vhd:1639:73  */
  assign n1543 = ea_register == 3'b100;
  assign n1544 = {n1543, n1540, n1538, n1536, n1534};
  /* TG68K_FPU.vhd:1624:65  */
  always @*
    case (n1544)
      5'b10000: n1547 = movem_predecrement;
      5'b01000: n1547 = movem_predecrement;
      5'b00100: n1547 = movem_predecrement;
      5'b00010: n1547 = 1'b0;
      5'b00001: n1547 = 1'b0;
      default: n1547 = movem_predecrement;
    endcase
  /* TG68K_FPU.vhd:1624:65  */
  always @*
    case (n1544)
      5'b10000: n1550 = movem_postincrement;
      5'b01000: n1550 = movem_postincrement;
      5'b00100: n1550 = movem_postincrement;
      5'b00010: n1550 = 1'b0;
      5'b00001: n1550 = 1'b0;
      default: n1550 = movem_postincrement;
    endcase
  /* TG68K_FPU.vhd:1623:57  */
  assign n1552 = ea_mode == 3'b111;
  assign n1553 = {n1552, n1532, n1525, n1523, n1521, n1519};
  /* TG68K_FPU.vhd:1598:57  */
  always @*
    case (n1553)
      6'b100000: n1559 = n1547;
      6'b010000: n1559 = 1'b0;
      6'b001000: n1559 = 1'b0;
      6'b000100: n1559 = 1'b1;
      6'b000010: n1559 = 1'b0;
      6'b000001: n1559 = 1'b0;
      default: n1559 = movem_predecrement;
    endcase
  /* TG68K_FPU.vhd:1598:57  */
  always @*
    case (n1553)
      6'b100000: n1565 = n1550;
      6'b010000: n1565 = 1'b0;
      6'b001000: n1565 = 1'b0;
      6'b000100: n1565 = 1'b0;
      6'b000010: n1565 = 1'b1;
      6'b000001: n1565 = 1'b0;
      default: n1565 = movem_postincrement;
    endcase
  /* TG68K_FPU.vhd:1657:57  */
  assign n1567 = movem_unit_address_error ? 1'b1 : n910;
  /* TG68K_FPU.vhd:1657:57  */
  assign n1570 = movem_unit_address_error ? 4'b1000 : 4'b1011;
  /* TG68K_FPU.vhd:1657:57  */
  assign n1572 = movem_unit_address_error ? 8'b00000011 : n913;
  /* TG68K_FPU.vhd:1585:49  */
  assign n1574 = n1515 ? 1'b1 : n1567;
  /* TG68K_FPU.vhd:1585:49  */
  assign n1576 = n1515 ? 4'b1000 : n1570;
  /* TG68K_FPU.vhd:1585:49  */
  assign n1577 = n1515 ? movem_register_list : n1516;
  /* TG68K_FPU.vhd:1585:49  */
  assign n1578 = n1515 ? movem_direction : n1517;
  /* TG68K_FPU.vhd:1585:49  */
  assign n1580 = n1515 ? 8'b00001100 : n1572;
  /* TG68K_FPU.vhd:1585:49  */
  assign n1581 = n1515 ? movem_predecrement : n1559;
  /* TG68K_FPU.vhd:1585:49  */
  assign n1582 = n1515 ? movem_postincrement : n1565;
  /* TG68K_FPU.vhd:1666:72  */
  assign n1584 = decoder_instruction_type == 4'b1001;
  /* TG68K_FPU.vhd:1683:72  */
  assign n1589 = decoder_instruction_type == 4'b0110;
  /* TG68K_FPU.vhd:1685:76  */
  assign n1590 = ~supervisor_mode;
  /* TG68K_FPU.vhd:1699:100  */
  assign n1592 = {fsave_frame_format, 24'b000000000000000000000000};
  /* TG68K_FPU.vhd:1685:57  */
  assign n1594 = n1590 ? 32'b00000000000000000000000000000000 : n1592;
  /* TG68K_FPU.vhd:1685:57  */
  assign n1596 = n1590 ? 1'b1 : n910;
  /* TG68K_FPU.vhd:1685:57  */
  assign n1599 = n1590 ? 4'b1000 : 4'b1001;
  /* TG68K_FPU.vhd:1685:57  */
  assign n1601 = n1590 ? fsave_frame_format_latched : fsave_frame_format;
  /* TG68K_FPU.vhd:1685:57  */
  assign n1603 = n1590 ? fsave_counter : 6'b000000;
  /* TG68K_FPU.vhd:1685:57  */
  assign n1605 = n1590 ? 8'b00100000 : n913;
  /* TG68K_FPU.vhd:1702:80  */
  assign n1607 = decoder_instruction_type == 4'b0111;
  /* TG68K_FPU.vhd:1704:76  */
  assign n1608 = ~supervisor_mode;
  /* TG68K_FPU.vhd:1704:57  */
  assign n1610 = n1608 ? 1'b1 : n910;
  /* TG68K_FPU.vhd:1704:57  */
  assign n1613 = n1608 ? 4'b1000 : 4'b1010;
  /* TG68K_FPU.vhd:1704:57  */
  assign n1615 = n1608 ? fsave_counter : 6'b000000;
  /* TG68K_FPU.vhd:1704:57  */
  assign n1617 = n1608 ? frestore_frame_format : 8'b00000000;
  /* TG68K_FPU.vhd:1704:57  */
  assign n1623 = n1608 ? 8'b00100000 : n913;
  /* TG68K_FPU.vhd:1718:80  */
  assign n1625 = decoder_instruction_type == 4'b0011;
  /* TG68K_FPU.vhd:1728:67  */
  assign n1626 = opcode[5:3]; // extract
  /* TG68K_FPU.vhd:1728:80  */
  assign n1628 = n1626 == 3'b010;
  /* TG68K_FPU.vhd:1728:98  */
  assign n1629 = opcode[2:0]; // extract
  /* TG68K_FPU.vhd:1728:111  */
  assign n1631 = n1629 == 3'b101;
  /* TG68K_FPU.vhd:1728:88  */
  assign n1632 = n1631 & n1628;
  /* TG68K_FPU.vhd:1730:83  */
  assign n1634 = extension_word == 16'b1110000011111111;
  /* TG68K_FPU.vhd:1735:86  */
  assign n1636 = extension_word == 16'b1011110000000000;
  /* TG68K_FPU.vhd:1737:92  */
  assign n1637 = ~supervisor_mode;
  /* TG68K_FPU.vhd:1735:65  */
  assign n1639 = n1650 ? 1'b1 : n910;
  /* TG68K_FPU.vhd:1737:73  */
  assign n1642 = n1637 ? 4'b1000 : 4'b1100;
  /* TG68K_FPU.vhd:1737:73  */
  assign n1644 = n1637 ? movem_direction : 1'b0;
  /* TG68K_FPU.vhd:1735:65  */
  assign n1646 = n1654 ? 8'b00100000 : n913;
  /* TG68K_FPU.vhd:1735:65  */
  assign n1649 = n1636 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:1735:65  */
  assign n1650 = n1637 & n1636;
  /* TG68K_FPU.vhd:1735:65  */
  assign n1652 = n1636 ? n1642 : 4'b0000;
  /* TG68K_FPU.vhd:1735:65  */
  assign n1653 = n1636 ? n1644 : movem_direction;
  /* TG68K_FPU.vhd:1735:65  */
  assign n1654 = n1637 & n1636;
  /* TG68K_FPU.vhd:1730:65  */
  assign n1656 = n1634 ? 1'b0 : n1649;
  /* TG68K_FPU.vhd:1730:65  */
  assign n1657 = n1634 ? n910 : n1639;
  /* TG68K_FPU.vhd:1730:65  */
  assign n1659 = n1634 ? 4'b1011 : n1652;
  /* TG68K_FPU.vhd:1730:65  */
  assign n1661 = n1634 ? 8'b11111111 : movem_register_list;
  /* TG68K_FPU.vhd:1730:65  */
  assign n1663 = n1634 ? 1'b0 : n1653;
  /* TG68K_FPU.vhd:1730:65  */
  assign n1664 = n1634 ? n913 : n1646;
  /* TG68K_FPU.vhd:1752:70  */
  assign n1665 = opcode[5:3]; // extract
  /* TG68K_FPU.vhd:1752:83  */
  assign n1667 = n1665 == 3'b001;
  /* TG68K_FPU.vhd:1752:101  */
  assign n1668 = opcode[2:0]; // extract
  /* TG68K_FPU.vhd:1752:114  */
  assign n1670 = n1668 == 3'b101;
  /* TG68K_FPU.vhd:1752:91  */
  assign n1671 = n1670 & n1667;
  /* TG68K_FPU.vhd:1754:83  */
  assign n1673 = extension_word == 16'b1101000011111111;
  /* TG68K_FPU.vhd:1759:86  */
  assign n1675 = extension_word == 16'b1001110000000000;
  /* TG68K_FPU.vhd:1761:92  */
  assign n1676 = ~supervisor_mode;
  /* TG68K_FPU.vhd:1759:65  */
  assign n1678 = n1689 ? 1'b1 : n910;
  /* TG68K_FPU.vhd:1761:73  */
  assign n1681 = n1676 ? 4'b1000 : 4'b1100;
  /* TG68K_FPU.vhd:1761:73  */
  assign n1683 = n1676 ? movem_direction : 1'b1;
  /* TG68K_FPU.vhd:1759:65  */
  assign n1685 = n1693 ? 8'b00100000 : n913;
  /* TG68K_FPU.vhd:1759:65  */
  assign n1688 = n1675 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:1759:65  */
  assign n1689 = n1676 & n1675;
  /* TG68K_FPU.vhd:1759:65  */
  assign n1691 = n1675 ? n1681 : 4'b0000;
  /* TG68K_FPU.vhd:1759:65  */
  assign n1692 = n1675 ? n1683 : movem_direction;
  /* TG68K_FPU.vhd:1759:65  */
  assign n1693 = n1676 & n1675;
  /* TG68K_FPU.vhd:1754:65  */
  assign n1695 = n1673 ? 1'b0 : n1688;
  /* TG68K_FPU.vhd:1754:65  */
  assign n1696 = n1673 ? n910 : n1678;
  /* TG68K_FPU.vhd:1754:65  */
  assign n1698 = n1673 ? 4'b1011 : n1691;
  /* TG68K_FPU.vhd:1752:57  */
  assign n1700 = n1709 ? 8'b11111111 : movem_register_list;
  /* TG68K_FPU.vhd:1754:65  */
  assign n1702 = n1673 ? 1'b1 : n1692;
  /* TG68K_FPU.vhd:1754:65  */
  assign n1703 = n1673 ? n913 : n1685;
  /* TG68K_FPU.vhd:1752:57  */
  assign n1705 = n1671 ? n1695 : 1'b1;
  /* TG68K_FPU.vhd:1752:57  */
  assign n1706 = n1671 ? n1696 : n910;
  /* TG68K_FPU.vhd:1752:57  */
  assign n1708 = n1671 ? n1698 : 4'b0000;
  /* TG68K_FPU.vhd:1752:57  */
  assign n1709 = n1673 & n1671;
  /* TG68K_FPU.vhd:1752:57  */
  assign n1710 = n1671 ? n1702 : movem_direction;
  /* TG68K_FPU.vhd:1752:57  */
  assign n1711 = n1671 ? n1703 : n913;
  /* TG68K_FPU.vhd:1728:57  */
  assign n1712 = n1632 ? n1656 : n1705;
  /* TG68K_FPU.vhd:1728:57  */
  assign n1713 = n1632 ? n1657 : n1706;
  /* TG68K_FPU.vhd:1728:57  */
  assign n1714 = n1632 ? n1659 : n1708;
  /* TG68K_FPU.vhd:1728:57  */
  assign n1715 = n1632 ? n1661 : n1700;
  /* TG68K_FPU.vhd:1728:57  */
  assign n1716 = n1632 ? n1663 : n1710;
  /* TG68K_FPU.vhd:1728:57  */
  assign n1717 = n1632 ? n1664 : n1711;
  /* TG68K_FPU.vhd:1780:80  */
  assign n1719 = decoder_instruction_type == 4'b0100;
  /* TG68K_FPU.vhd:1782:74  */
  assign n1720 = extension_word[15:13]; // extract
  /* TG68K_FPU.vhd:1782:89  */
  assign n1722 = n1720 == 3'b100;
  /* TG68K_FPU.vhd:1784:82  */
  assign n1723 = extension_word[13]; // extract
  /* TG68K_FPU.vhd:1784:87  */
  assign n1724 = ~n1723;
  /* TG68K_FPU.vhd:1786:92  */
  assign n1725 = extension_word[12:10]; // extract
  /* TG68K_FPU.vhd:1787:81  */
  assign n1727 = n1725 == 3'b001;
  /* TG68K_FPU.vhd:1789:81  */
  assign n1729 = n1725 == 3'b010;
  /* TG68K_FPU.vhd:1791:81  */
  assign n1731 = n1725 == 3'b100;
  assign n1732 = {n1731, n1729, n1727};
  /* TG68K_FPU.vhd:1786:73  */
  always @*
    case (n1732)
      3'b100: n1734 = fpiar;
      3'b010: n1734 = fpsr;
      3'b001: n1734 = fpcr;
      default: n1734 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:1800:92  */
  assign n1735 = extension_word[12:10]; // extract
  /* TG68K_FPU.vhd:597:30  */
  assign n1743 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:43  */
  assign n1745 = n1743 == 2'b11;
  assign n1747 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:17  */
  assign n1748 = n1745 ? 2'b00 : n1747;
  assign n1752 = cpu_data_in[15:8]; // extract
  assign n1754 = {16'b0000000000000000, n1752, n1748, 6'b000000};
  /* TG68K_FPU.vhd:1801:81  */
  assign n1756 = n1735 == 3'b001;
  /* TG68K_FPU.vhd:1803:81  */
  assign n1765 = n1735 == 3'b010;
  /* TG68K_FPU.vhd:1805:81  */
  assign n1767 = n1735 == 3'b100;
  assign n1768 = {n1767, n1765, n1756};
  /* TG68K_FPU.vhd:1800:73  */
  always @*
    case (n1768)
      3'b100: n1769 = fpcr;
      3'b010: n1769 = fpcr;
      3'b001: n1769 = n1754;
      default: n1769 = fpcr;
    endcase
  /* TG68K_FPU.vhd:1800:73  */
  always @*
    case (n1768)
      3'b100: n1770 = fpsr;
      3'b010: n1770 = cpu_data_in;
      3'b001: n1770 = fpsr;
      default: n1770 = fpsr;
    endcase
  /* TG68K_FPU.vhd:1800:73  */
  always @*
    case (n1768)
      3'b100: n1771 = cpu_data_in;
      3'b010: n1771 = n919;
      3'b001: n1771 = n919;
      default: n1771 = n919;
    endcase
  /* TG68K_FPU.vhd:1784:65  */
  assign n1773 = n1724 ? n1734 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1784:65  */
  assign n1774 = n1724 ? fpcr : n1769;
  /* TG68K_FPU.vhd:1784:65  */
  assign n1775 = n1724 ? fpsr : n1770;
  /* TG68K_FPU.vhd:1784:65  */
  assign n1776 = n1724 ? n919 : n1771;
  /* TG68K_FPU.vhd:1782:57  */
  assign n1778 = n1722 ? n1773 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1780:49  */
  assign n1779 = n2289 ? n1774 : fpcr;
  /* TG68K_FPU.vhd:1780:49  */
  assign n1780 = n2290 ? n1775 : fpsr;
  /* TG68K_FPU.vhd:1780:49  */
  assign n1781 = n2291 ? n1776 : n919;
  /* TG68K_FPU.vhd:1818:80  */
  assign n1783 = decoder_instruction_type == 4'b0000;
  /* TG68K_FPU.vhd:1821:74  */
  assign n1785 = fpu_operation == 7'b0000000;
  /* TG68K_FPU.vhd:1821:102  */
  assign n1787 = fpu_operation == 7'b0000001;
  /* TG68K_FPU.vhd:1821:85  */
  assign n1788 = n1785 | n1787;
  /* TG68K_FPU.vhd:1821:129  */
  assign n1790 = fpu_operation == 7'b0000011;
  /* TG68K_FPU.vhd:1821:112  */
  assign n1791 = n1788 | n1790;
  /* TG68K_FPU.vhd:1822:69  */
  assign n1793 = fpu_operation == 7'b0100010;
  /* TG68K_FPU.vhd:1821:141  */
  assign n1794 = n1791 | n1793;
  /* TG68K_FPU.vhd:1822:96  */
  assign n1796 = fpu_operation == 7'b0101000;
  /* TG68K_FPU.vhd:1822:79  */
  assign n1797 = n1794 | n1796;
  /* TG68K_FPU.vhd:1822:123  */
  assign n1799 = fpu_operation == 7'b0100011;
  /* TG68K_FPU.vhd:1822:106  */
  assign n1800 = n1797 | n1799;
  /* TG68K_FPU.vhd:1823:69  */
  assign n1802 = fpu_operation == 7'b0100000;
  /* TG68K_FPU.vhd:1822:133  */
  assign n1803 = n1800 | n1802;
  /* TG68K_FPU.vhd:1823:96  */
  assign n1805 = fpu_operation == 7'b0000100;
  /* TG68K_FPU.vhd:1823:79  */
  assign n1806 = n1803 | n1805;
  /* TG68K_FPU.vhd:1824:69  */
  assign n1808 = fpu_operation == 7'b0011000;
  /* TG68K_FPU.vhd:1823:107  */
  assign n1809 = n1806 | n1808;
  /* TG68K_FPU.vhd:1824:96  */
  assign n1811 = fpu_operation == 7'b0011010;
  /* TG68K_FPU.vhd:1824:79  */
  assign n1812 = n1809 | n1811;
  /* TG68K_FPU.vhd:1825:69  */
  assign n1814 = fpu_operation == 7'b0111000;
  /* TG68K_FPU.vhd:1824:106  */
  assign n1815 = n1812 | n1814;
  /* TG68K_FPU.vhd:1825:96  */
  assign n1817 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:1825:79  */
  assign n1818 = n1815 | n1817;
  /* TG68K_FPU.vhd:1826:69  */
  assign n1820 = fpu_operation == 7'b0100100;
  /* TG68K_FPU.vhd:1825:106  */
  assign n1821 = n1818 | n1820;
  /* TG68K_FPU.vhd:1826:99  */
  assign n1823 = fpu_operation == 7'b0100111;
  /* TG68K_FPU.vhd:1826:82  */
  assign n1824 = n1821 | n1823;
  /* TG68K_FPU.vhd:1827:69  */
  assign n1826 = fpu_operation == 7'b0001110;
  /* TG68K_FPU.vhd:1826:112  */
  assign n1827 = n1824 | n1826;
  /* TG68K_FPU.vhd:1827:96  */
  assign n1829 = fpu_operation == 7'b0011101;
  /* TG68K_FPU.vhd:1827:79  */
  assign n1830 = n1827 | n1829;
  /* TG68K_FPU.vhd:1827:123  */
  assign n1832 = fpu_operation == 7'b0001111;
  /* TG68K_FPU.vhd:1827:106  */
  assign n1833 = n1830 | n1832;
  /* TG68K_FPU.vhd:1828:69  */
  assign n1835 = fpu_operation == 7'b0001100;
  /* TG68K_FPU.vhd:1827:133  */
  assign n1836 = n1833 | n1835;
  /* TG68K_FPU.vhd:1828:97  */
  assign n1838 = fpu_operation == 7'b0011100;
  /* TG68K_FPU.vhd:1828:80  */
  assign n1839 = n1836 | n1838;
  /* TG68K_FPU.vhd:1828:125  */
  assign n1841 = fpu_operation == 7'b0001010;
  /* TG68K_FPU.vhd:1828:108  */
  assign n1842 = n1839 | n1841;
  /* TG68K_FPU.vhd:1829:69  */
  assign n1844 = fpu_operation == 7'b0001011;
  /* TG68K_FPU.vhd:1828:136  */
  assign n1845 = n1842 | n1844;
  /* TG68K_FPU.vhd:1829:97  */
  assign n1847 = fpu_operation == 7'b0011001;
  /* TG68K_FPU.vhd:1829:80  */
  assign n1848 = n1845 | n1847;
  /* TG68K_FPU.vhd:1829:125  */
  assign n1850 = fpu_operation == 7'b0001001;
  /* TG68K_FPU.vhd:1829:108  */
  assign n1851 = n1848 | n1850;
  /* TG68K_FPU.vhd:1830:69  */
  assign n1853 = fpu_operation == 7'b0001101;
  /* TG68K_FPU.vhd:1829:136  */
  assign n1854 = n1851 | n1853;
  /* TG68K_FPU.vhd:1830:98  */
  assign n1856 = fpu_operation == 7'b0010000;
  /* TG68K_FPU.vhd:1830:81  */
  assign n1857 = n1854 | n1856;
  /* TG68K_FPU.vhd:1830:126  */
  assign n1859 = fpu_operation == 7'b0000111;
  /* TG68K_FPU.vhd:1830:109  */
  assign n1860 = n1857 | n1859;
  /* TG68K_FPU.vhd:1831:69  */
  assign n1862 = fpu_operation == 7'b0010001;
  /* TG68K_FPU.vhd:1830:139  */
  assign n1863 = n1860 | n1862;
  /* TG68K_FPU.vhd:1831:99  */
  assign n1865 = fpu_operation == 7'b0010010;
  /* TG68K_FPU.vhd:1831:82  */
  assign n1866 = n1863 | n1865;
  /* TG68K_FPU.vhd:1831:129  */
  assign n1868 = fpu_operation == 7'b0010100;
  /* TG68K_FPU.vhd:1831:112  */
  assign n1869 = n1866 | n1868;
  /* TG68K_FPU.vhd:1832:69  */
  assign n1871 = fpu_operation == 7'b0000101;
  /* TG68K_FPU.vhd:1831:140  */
  assign n1872 = n1869 | n1871;
  /* TG68K_FPU.vhd:1832:99  */
  assign n1874 = fpu_operation == 7'b0010101;
  /* TG68K_FPU.vhd:1832:82  */
  assign n1875 = n1872 | n1874;
  /* TG68K_FPU.vhd:1833:69  */
  assign n1877 = fpu_operation == 7'b0010110;
  /* TG68K_FPU.vhd:1832:111  */
  assign n1878 = n1875 | n1877;
  /* TG68K_FPU.vhd:1833:97  */
  assign n1880 = fpu_operation == 7'b1000001;
  /* TG68K_FPU.vhd:1833:80  */
  assign n1881 = n1878 | n1880;
  /* TG68K_FPU.vhd:1833:127  */
  assign n1883 = fpu_operation == 7'b0100001;
  /* TG68K_FPU.vhd:1833:110  */
  assign n1884 = n1881 | n1883;
  /* TG68K_FPU.vhd:1834:69  */
  assign n1886 = fpu_operation == 7'b0100101;
  /* TG68K_FPU.vhd:1833:137  */
  assign n1887 = n1884 | n1886;
  /* TG68K_FPU.vhd:1834:96  */
  assign n1889 = fpu_operation == 7'b0100110;
  /* TG68K_FPU.vhd:1834:79  */
  assign n1890 = n1887 | n1889;
  /* TG68K_FPU.vhd:1834:125  */
  assign n1892 = fpu_operation == 7'b0011110;
  /* TG68K_FPU.vhd:1834:108  */
  assign n1893 = n1890 | n1892;
  /* TG68K_FPU.vhd:1835:69  */
  assign n1895 = fpu_operation == 7'b0011111;
  /* TG68K_FPU.vhd:1834:138  */
  assign n1896 = n1893 | n1895;
  /* TG68K_FPU.vhd:1835:99  */
  assign n1898 = fpu_operation == 7'b0110000;
  /* TG68K_FPU.vhd:1835:82  */
  assign n1899 = n1896 | n1898;
  /* TG68K_FPU.vhd:1856:82  */
  assign n1927 = fpu_operation == 7'b1000001;
  /* TG68K_FPU.vhd:1858:101  */
  assign n1928 = extension_word[6:0]; // extract
  /* TG68K_FPU.vhd:1861:85  */
  assign n1930 = fpu_operation == 7'b0000010;
  /* TG68K_FPU.vhd:1866:85  */
  assign n1932 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:1866:112  */
  assign n1934 = fpu_operation == 7'b0111000;
  /* TG68K_FPU.vhd:1866:95  */
  assign n1935 = n1932 | n1934;
  /* TG68K_FPU.vhd:1869:108  */
  assign n1937 = cir_address == 5'b00101;
  /* TG68K_FPU.vhd:1869:92  */
  assign n1938 = n1937 & cir_write;
  /* TG68K_FPU.vhd:1869:73  */
  assign n1941 = n1938 ? 4'b0101 : 4'b0010;
  /* TG68K_FPU.vhd:1866:65  */
  assign n1943 = n1935 ? n1941 : 4'b0010;
  /* TG68K_FPU.vhd:1861:65  */
  assign n1946 = n1930 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:1861:65  */
  assign n1948 = n1930 ? 4'b0000 : n1943;
  /* TG68K_FPU.vhd:1856:65  */
  assign n1950 = n1927 ? 1'b0 : n1946;
  /* TG68K_FPU.vhd:1856:65  */
  assign n1952 = n1927 ? 4'b0110 : n1948;
  /* TG68K_FPU.vhd:1818:49  */
  assign n1953 = n2278 ? n1928 : rom_offset;
  /* TG68K_FPU.vhd:1818:49  */
  assign n1955 = n2279 ? 1'b1 : rom_read_enable;
  /* TG68K_FPU.vhd:1821:57  */
  assign n1957 = n1899 ? n1950 : 1'b0;
  /* TG68K_FPU.vhd:1821:57  */
  assign n1959 = n1899 ? n910 : 1'b1;
  /* TG68K_FPU.vhd:1821:57  */
  assign n1961 = n1899 ? n1952 : 4'b1000;
  /* TG68K_FPU.vhd:1821:57  */
  assign n1963 = n1899 ? n913 : 8'b00001100;
  /* TG68K_FPU.vhd:1821:57  */
  assign n1964 = n1927 & n1899;
  /* TG68K_FPU.vhd:1821:57  */
  assign n1965 = n1927 & n1899;
  /* TG68K_FPU.vhd:1886:80  */
  assign n1967 = decoder_instruction_type == 4'b0001;
  /* TG68K_FPU.vhd:1891:60  */
  assign n1968 = {28'b0, decoder_source_reg};  //  uext
  /* TG68K_FPU.vhd:1891:101  */
  assign n1969 = {1'b0, n1968};  //  uext
  /* TG68K_FPU.vhd:1891:101  */
  assign n1971 = $signed(n1969) > $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:1891:57  */
  assign n1973 = n1971 ? 1'b1 : n910;
  /* TG68K_FPU.vhd:1891:57  */
  assign n1977 = n1971 ? 8'b00001100 : n913;
  /* TG68K_FPU.vhd:1905:102  */
  assign n1980 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1906:118  */
  assign n1985 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1906:159  */
  assign n1987 = fp_registers[n6897 + 65 +: 7]; //(dyn_extract)
  /* TG68K_FPU.vhd:1905:148  */
  assign n1988 = {n6894, n1987};
  /* TG68K_FPU.vhd:1906:174  */
  assign n1990 = {n1988, 1'b1};
  /* TG68K_FPU.vhd:1907:118  */
  assign n1993 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1907:159  */
  assign n1995 = fp_registers[n6900 + 41 +: 23]; //(dyn_extract)
  /* TG68K_FPU.vhd:1906:180  */
  assign n1996 = {n1990, n1995};
  /* TG68K_FPU.vhd:1898:65  */
  assign n1998 = decoder_dest_format == 3'b001;
  /* TG68K_FPU.vhd:1916:102  */
  assign n2001 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1917:118  */
  assign n2006 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1916:148  */
  assign n2009 = {n6905, n6910};
  /* TG68K_FPU.vhd:1917:174  */
  assign n2011 = {n2009, 1'b0};
  /* TG68K_FPU.vhd:1918:118  */
  assign n2014 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1917:180  */
  assign n2017 = {n2011, n6915};
  /* TG68K_FPU.vhd:1909:65  */
  assign n2019 = decoder_dest_format == 3'b101;
  /* TG68K_FPU.vhd:1933:89  */
  assign n2037 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1933:130  */
  assign n2039 = fp_registers[n6918 + 64 +: 15]; //(dyn_extract)
  /* TG68K_FPU.vhd:1933:145  */
  assign n2041 = n2039 == 15'b000000000000000;
  /* TG68K_FPU.vhd:1936:92  */
  assign n2044 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1936:133  */
  assign n2046 = fp_registers[n6921 + 64 +: 15]; //(dyn_extract)
  /* TG68K_FPU.vhd:1936:148  */
  assign n2048 = n2046 == 15'b111111111111111;
  /* TG68K_FPU.vhd:1938:97  */
  assign n2051 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1938:81  */
  assign n2056 = n6926 ? 32'b10000000000000000000000000000000 : 32'b01111111111111111111111111111111;
  /* TG68K_FPU.vhd:1947:117  */
  assign n2059 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1947:158  */
  assign n2061 = fp_registers[n6929 + 64 +: 15]; //(dyn_extract)
  /* TG68K_FPU.vhd:1947:84  */
  assign n2062 = {16'b0, n2061};  //  uext
  /* TG68K_FPU.vhd:1947:175  */
  assign n2063 = {1'b0, n2062};  //  uext
  /* TG68K_FPU.vhd:1947:175  */
  assign n2065 = $signed(n2063) < $signed(32'b00000000000000000011111111111111);
  /* TG68K_FPU.vhd:1950:120  */
  assign n2068 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1950:161  */
  assign n2070 = fp_registers[n6932 + 64 +: 15]; //(dyn_extract)
  /* TG68K_FPU.vhd:1950:87  */
  assign n2071 = {16'b0, n2070};  //  uext
  /* TG68K_FPU.vhd:1950:178  */
  assign n2072 = {1'b0, n2071};  //  uext
  /* TG68K_FPU.vhd:1950:178  */
  assign n2074 = $signed(n2072) > $signed(32'b00000000000000000100000000011101);
  /* TG68K_FPU.vhd:1952:105  */
  assign n2077 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1952:89  */
  assign n2082 = n6937 ? 32'b10000000000000000000000000000000 : 32'b01111111111111111111111111111111;
  /* TG68K_FPU.vhd:1960:125  */
  assign n2085 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1960:166  */
  assign n2087 = fp_registers[n6940 + 64 +: 15]; //(dyn_extract)
  /* TG68K_FPU.vhd:1960:92  */
  assign n2088 = {16'b0, n2087};  //  uext
  /* TG68K_FPU.vhd:1960:183  */
  assign n2089 = {1'b0, n2088};  //  uext
  /* TG68K_FPU.vhd:1960:183  */
  assign n2091 = $signed(n2089) < $signed(32'b00000000000000000011111111100000);
  /* TG68K_FPU.vhd:1963:128  */
  assign n2094 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1963:169  */
  assign n2096 = fp_registers[n6943 + 64 +: 15]; //(dyn_extract)
  /* TG68K_FPU.vhd:1963:95  */
  assign n2097 = {16'b0, n2096};  //  uext
  /* TG68K_FPU.vhd:1963:186  */
  assign n2098 = {1'b0, n2097};  //  uext
  /* TG68K_FPU.vhd:1963:186  */
  assign n2100 = $signed(n2098) > $signed(32'b00000000000000000100000000011101);
  /* TG68K_FPU.vhd:1968:155  */
  assign n2103 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1968:196  */
  assign n2105 = fp_registers[n6946 + 64 +: 15]; //(dyn_extract)
  /* TG68K_FPU.vhd:1968:122  */
  assign n2106 = {16'b0, n2105};  //  uext
  /* TG68K_FPU.vhd:1968:213  */
  assign n2107 = {1'b0, n2106};  //  uext
  /* TG68K_FPU.vhd:1968:213  */
  assign n2109 = n2107 - 32'b00000000000000000011111111111111;
  /* TG68K_FPU.vhd:1968:119  */
  assign n2111 = 32'b00000000000000000000000000111111 - n2109;
  /* TG68K_FPU.vhd:1968:116  */
  assign n2112 = n2111[5:0];  // trunc
  /* TG68K_FPU.vhd:1963:89  */
  assign n2114 = n2100 ? 6'b000000 : n2112;
  /* TG68K_FPU.vhd:1960:89  */
  assign n2116 = n2091 ? 6'b111111 : n2114;
  /* TG68K_FPU.vhd:1974:108  */
  assign n2117 = {26'b0, fp_to_int_shift};  //  uext
  /* TG68K_FPU.vhd:1974:108  */
  assign n2119 = $signed(n2117) <= $signed(32'b00000000000000000000000000011111);
  /* TG68K_FPU.vhd:1978:146  */
  assign n2122 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1978:187  */
  assign n2124 = fp_registers[n6949 + 32 +: 32]; //(dyn_extract)
  /* TG68K_FPU.vhd:1977:105  */
  assign n2126 = fp_to_int_shift == 6'b000000;
  /* TG68K_FPU.vhd:1981:184  */
  assign n2129 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1981:225  */
  assign n2131 = fp_registers[n6952 + 0 +: 64]; //(dyn_extract)
  /* TG68K_FPU.vhd:1981:241  */
  assign n2132 = {25'b0, fp_to_int_shift};  //  uext
  /* TG68K_FPU.vhd:1981:150  */
  assign n2133 = n2131 >> n2132;
  /* TG68K_FPU.vhd:1981:257  */
  assign n2134 = n2133[31:0]; // extract
  /* TG68K_FPU.vhd:1979:105  */
  assign n2137 = $unsigned(fp_to_int_shift) >= $unsigned(6'b000001);
  /* TG68K_FPU.vhd:1979:105  */
  assign n2138 = $unsigned(fp_to_int_shift) <= $unsigned(6'b011111);
  /* TG68K_FPU.vhd:1979:105  */
  assign n2139 = n2137 & n2138;
  assign n2140 = {n2139, n2126};
  /* TG68K_FPU.vhd:1976:97  */
  always @*
    case (n2140)
      2'b10: n2142 = n2134;
      2'b01: n2142 = n2124;
      default: n2142 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:1974:89  */
  assign n2144 = n2119 ? n2142 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1991:105  */
  assign n2147 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:1992:139  */
  assign n2150 = ~fp_to_int_result;
  /* TG68K_FPU.vhd:1992:161  */
  assign n2152 = n2150 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:1991:89  */
  assign n2153 = n6957 ? n2152 : fp_to_int_result;
  /* TG68K_FPU.vhd:1950:81  */
  assign n2154 = n2074 ? n2082 : n2153;
  /* TG68K_FPU.vhd:1950:81  */
  assign n2155 = n2074 ? fp_to_int_shift : n2116;
  /* TG68K_FPU.vhd:1950:81  */
  assign n2156 = n2074 ? fp_to_int_result : n2144;
  /* TG68K_FPU.vhd:1947:81  */
  assign n2158 = n2065 ? 32'b00000000000000000000000000000000 : n2154;
  /* TG68K_FPU.vhd:1947:81  */
  assign n2159 = n2065 ? fp_to_int_shift : n2155;
  /* TG68K_FPU.vhd:1947:81  */
  assign n2160 = n2065 ? fp_to_int_result : n2156;
  /* TG68K_FPU.vhd:1936:73  */
  assign n2161 = n2048 ? n2056 : n2158;
  /* TG68K_FPU.vhd:1936:73  */
  assign n2162 = n2048 ? fp_to_int_shift : n2159;
  /* TG68K_FPU.vhd:1936:73  */
  assign n2163 = n2048 ? fp_to_int_result : n2160;
  /* TG68K_FPU.vhd:1933:73  */
  assign n2165 = n2041 ? 32'b00000000000000000000000000000000 : n2161;
  /* TG68K_FPU.vhd:1933:73  */
  assign n2166 = n2041 ? fp_to_int_shift : n2162;
  /* TG68K_FPU.vhd:1933:73  */
  assign n2167 = n2041 ? fp_to_int_result : n2163;
  /* TG68K_FPU.vhd:1920:65  */
  assign n2169 = decoder_dest_format == 3'b000;
  /* TG68K_FPU.vhd:2006:120  */
  assign n2172 = 3'b111 - decoder_source_reg;
  /* TG68K_FPU.vhd:2000:65  */
  assign n2177 = decoder_dest_format == 3'b011;
  /* TG68K_FPU.vhd:2014:120  */
  assign n2180 = 3'b111 - decoder_source_reg;
  assign n2184 = {n2177, n2169, n2019, n1998};
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2186 = 32'b00000000000000000000000000000000;
      4'b0100: n2186 = n2165;
      4'b0010: n2186 = n2017;
      4'b0001: n2186 = n1996;
      default: n2186 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2189 = 1'b1;
      4'b0100: n2189 = converter_start;
      4'b0010: n2189 = converter_start;
      4'b0001: n2189 = converter_start;
      default: n2189 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2192 = 3'b010;
      4'b0100: n2192 = converter_source_format;
      4'b0010: n2192 = converter_source_format;
      4'b0001: n2192 = converter_source_format;
      default: n2192 = 3'b010;
    endcase
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2195 = 3'b011;
      4'b0100: n2195 = converter_dest_format;
      4'b0010: n2195 = converter_dest_format;
      4'b0001: n2195 = converter_dest_format;
      default: n2195 = 3'b010;
    endcase
  assign n2196 = converter_data_in[79:0]; // extract
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2197 = n6958;
      4'b0100: n2197 = n2196;
      4'b0010: n2197 = n2196;
      4'b0001: n2197 = n2196;
      default: n2197 = n6959;
    endcase
  assign n2198 = converter_data_in[95:80]; // extract
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2199 = 16'b0000000000000000;
      4'b0100: n2199 = n2198;
      4'b0010: n2199 = n2198;
      4'b0001: n2199 = n2198;
      default: n2199 = 16'b0000000000000000;
    endcase
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2203 = fp_to_int_shift;
      4'b0100: n2203 = n2166;
      4'b0010: n2203 = fp_to_int_shift;
      4'b0001: n2203 = fp_to_int_shift;
      default: n2203 = fp_to_int_shift;
    endcase
  /* TG68K_FPU.vhd:1897:57  */
  always @*
    case (n2184)
      4'b1000: n2204 = fp_to_int_result;
      4'b0100: n2204 = n2167;
      4'b0010: n2204 = fp_to_int_result;
      4'b0001: n2204 = fp_to_int_result;
      default: n2204 = fp_to_int_result;
    endcase
  /* TG68K_FPU.vhd:2019:80  */
  assign n2206 = decoder_instruction_type == 4'b0010;
  /* TG68K_FPU.vhd:2023:65  */
  assign n2208 = decoder_source_format == 3'b001;
  /* TG68K_FPU.vhd:2030:65  */
  assign n2210 = decoder_source_format == 3'b101;
  /* TG68K_FPU.vhd:2037:65  */
  assign n2212 = decoder_source_format == 3'b000;
  /* TG68K_FPU.vhd:2044:65  */
  assign n2214 = decoder_source_format == 3'b011;
  assign n2215 = {n2214, n2212, n2210, n2208};
  /* TG68K_FPU.vhd:2022:57  */
  always @*
    case (n2215)
      4'b1000: n2217 = converter_start;
      4'b0100: n2217 = converter_start;
      4'b0010: n2217 = converter_start;
      4'b0001: n2217 = converter_start;
      default: n2217 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:2022:57  */
  always @*
    case (n2215)
      4'b1000: n2219 = converter_source_format;
      4'b0100: n2219 = converter_source_format;
      4'b0010: n2219 = converter_source_format;
      4'b0001: n2219 = converter_source_format;
      default: n2219 = 3'b010;
    endcase
  /* TG68K_FPU.vhd:2022:57  */
  always @*
    case (n2215)
      4'b1000: n2221 = converter_dest_format;
      4'b0100: n2221 = converter_dest_format;
      4'b0010: n2221 = converter_dest_format;
      4'b0001: n2221 = converter_dest_format;
      default: n2221 = 3'b010;
    endcase
  /* TG68K_FPU.vhd:2064:80  */
  assign n2223 = decoder_instruction_type == 4'b0011;
  /* TG68K_FPU.vhd:2069:74  */
  assign n2224 = extension_word[7:0]; // extract
  /* TG68K_FPU.vhd:2069:87  */
  assign n2226 = n2224 == 8'b00000000;
  /* TG68K_FPU.vhd:2069:57  */
  assign n2229 = n2226 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:2069:57  */
  assign n2232 = n2226 ? 4'b0000 : 4'b0101;
  /* TG68K_FPU.vhd:2064:49  */
  assign n2234 = n2223 ? n2229 : 1'b0;
  /* TG68K_FPU.vhd:2064:49  */
  assign n2236 = n2223 ? n910 : 1'b1;
  /* TG68K_FPU.vhd:2064:49  */
  assign n2238 = n2223 ? n2232 : 4'b1000;
  /* TG68K_FPU.vhd:2064:49  */
  assign n2240 = n2223 ? n913 : 8'b00001100;
  /* TG68K_FPU.vhd:2019:49  */
  assign n2242 = n2206 ? 1'b0 : n2234;
  /* TG68K_FPU.vhd:2019:49  */
  assign n2243 = n2206 ? n910 : n2236;
  /* TG68K_FPU.vhd:2019:49  */
  assign n2245 = n2206 ? 4'b0011 : n2238;
  /* TG68K_FPU.vhd:2019:49  */
  assign n2246 = n2206 ? n913 : n2240;
  /* TG68K_FPU.vhd:2019:49  */
  assign n2247 = n2206 ? n2217 : converter_start;
  /* TG68K_FPU.vhd:2019:49  */
  assign n2248 = n2206 ? n2219 : converter_source_format;
  /* TG68K_FPU.vhd:2019:49  */
  assign n2249 = n2206 ? n2221 : converter_dest_format;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2251 = n1967 ? n2186 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2253 = n1967 ? 1'b0 : n2242;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2254 = n1967 ? n1973 : n2243;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2256 = n1967 ? 4'b0100 : n2245;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2257 = n1967 ? n1977 : n2246;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2258 = n1967 ? n2189 : n2247;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2259 = n1967 ? n2192 : n2248;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2260 = n1967 ? n2195 : n2249;
  assign n2261 = {n2199, n2197};
  /* TG68K_FPU.vhd:1886:49  */
  assign n2262 = n1967 ? n2261 : converter_data_in;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2266 = n1967 ? n2203 : fp_to_int_shift;
  /* TG68K_FPU.vhd:1886:49  */
  assign n2267 = n1967 ? n2204 : fp_to_int_result;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2269 = n1783 ? 32'b00000000000000000000000000000000 : n2251;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2270 = n1783 ? n1957 : n2253;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2271 = n1783 ? n1959 : n2254;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2272 = n1783 ? n1961 : n2256;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2273 = n1783 ? n1963 : n2257;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2274 = n1783 ? converter_start : n2258;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2275 = n1783 ? converter_source_format : n2259;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2276 = n1783 ? converter_dest_format : n2260;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2277 = n1783 ? converter_data_in : n2262;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2278 = n1964 & n1783;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2279 = n1965 & n1783;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2283 = n1783 ? fp_to_int_shift : n2266;
  /* TG68K_FPU.vhd:1818:49  */
  assign n2284 = n1783 ? fp_to_int_result : n2267;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2285 = n1719 ? n1778 : n2269;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2287 = n1719 ? 1'b1 : n2270;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2288 = n1719 ? n910 : n2271;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2289 = n1722 & n1719;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2290 = n1722 & n1719;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2291 = n1722 & n1719;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2293 = n1719 ? 4'b0000 : n2272;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2294 = n1719 ? n913 : n2273;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2295 = n1719 ? converter_start : n2274;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2296 = n1719 ? converter_source_format : n2275;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2297 = n1719 ? converter_dest_format : n2276;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2298 = n1719 ? converter_data_in : n2277;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2299 = n1719 ? rom_offset : n1953;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2300 = n1719 ? rom_read_enable : n1955;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2304 = n1719 ? fp_to_int_shift : n2283;
  /* TG68K_FPU.vhd:1780:49  */
  assign n2305 = n1719 ? fp_to_int_result : n2284;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2307 = n1625 ? 32'b00000000000000000000000000000000 : n2285;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2308 = n1625 ? n1712 : n2287;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2309 = n1625 ? n1713 : n2288;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2310 = n1625 ? fpcr : n1779;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2311 = n1625 ? fpsr : n1780;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2312 = n1625 ? n919 : n1781;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2313 = n1625 ? n1714 : n2293;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2314 = n1625 ? n1715 : movem_register_list;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2315 = n1625 ? n1716 : movem_direction;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2316 = n1625 ? n1717 : n2294;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2317 = n1625 ? converter_start : n2295;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2318 = n1625 ? converter_source_format : n2296;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2319 = n1625 ? converter_dest_format : n2297;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2320 = n1625 ? converter_data_in : n2298;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2321 = n1625 ? rom_offset : n2299;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2322 = n1625 ? rom_read_enable : n2300;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2326 = n1625 ? fp_to_int_shift : n2304;
  /* TG68K_FPU.vhd:1718:49  */
  assign n2327 = n1625 ? fp_to_int_result : n2305;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2329 = n1607 ? 32'b00000000000000000000000000000000 : n2307;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2331 = n1607 ? 1'b0 : n2308;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2332 = n1607 ? n1610 : n2309;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2333 = n1607 ? fpcr : n2310;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2334 = n1607 ? fpsr : n2311;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2335 = n1607 ? n919 : n2312;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2336 = n1607 ? n1613 : n2313;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2337 = n1607 ? movem_register_list : n2314;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2338 = n1607 ? movem_direction : n2315;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2339 = n1607 ? n1615 : fsave_counter;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2340 = n1607 ? n1617 : frestore_frame_format;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2343 = n1607 ? n1623 : n2316;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2344 = n1607 ? converter_start : n2317;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2345 = n1607 ? converter_source_format : n2318;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2346 = n1607 ? converter_dest_format : n2319;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2347 = n1607 ? converter_data_in : n2320;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2348 = n1607 ? rom_offset : n2321;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2349 = n1607 ? rom_read_enable : n2322;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2353 = n1607 ? fp_to_int_shift : n2326;
  /* TG68K_FPU.vhd:1702:49  */
  assign n2354 = n1607 ? fp_to_int_result : n2327;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2355 = n1589 ? n1594 : n2329;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2357 = n1589 ? 1'b0 : n2331;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2358 = n1589 ? n1596 : n2332;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2359 = n1589 ? fpcr : n2333;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2360 = n1589 ? fpsr : n2334;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2361 = n1589 ? n919 : n2335;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2362 = n1589 ? n1599 : n2336;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2364 = n1589 ? n1601 : fsave_frame_format_latched;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2365 = n1589 ? movem_register_list : n2337;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2366 = n1589 ? movem_direction : n2338;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2367 = n1589 ? n1603 : n2339;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2368 = n1589 ? frestore_frame_format : n2340;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2371 = n1589 ? n1605 : n2343;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2372 = n1589 ? converter_start : n2344;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2373 = n1589 ? converter_source_format : n2345;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2374 = n1589 ? converter_dest_format : n2346;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2375 = n1589 ? converter_data_in : n2347;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2376 = n1589 ? rom_offset : n2348;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2377 = n1589 ? rom_read_enable : n2349;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2381 = n1589 ? fp_to_int_shift : n2353;
  /* TG68K_FPU.vhd:1683:41  */
  assign n2382 = n1589 ? fp_to_int_result : n2354;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2384 = n1584 ? 32'b00000000000000000000000000000000 : n2355;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2386 = n1584 ? 1'b1 : n2357;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2387 = n1584 ? n910 : n2358;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2388 = n1584 ? fpcr : n2359;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2389 = n1584 ? fpsr : n2360;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2390 = n1584 ? n919 : n2361;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2392 = n1584 ? 4'b0000 : n2362;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2394 = n1584 ? fsave_frame_format_latched : n2364;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2395 = n1584 ? movem_register_list : n2365;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2396 = n1584 ? movem_direction : n2366;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2397 = n1584 ? fsave_counter : n2367;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2398 = n1584 ? frestore_frame_format : n2368;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2401 = n1584 ? n913 : n2371;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2402 = n1584 ? converter_start : n2372;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2403 = n1584 ? converter_source_format : n2373;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2404 = n1584 ? converter_dest_format : n2374;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2405 = n1584 ? converter_data_in : n2375;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2406 = n1584 ? rom_offset : n2376;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2407 = n1584 ? rom_read_enable : n2377;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2411 = n1584 ? fp_to_int_shift : n2381;
  /* TG68K_FPU.vhd:1666:41  */
  assign n2412 = n1584 ? fp_to_int_result : n2382;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2414 = n1500 ? 32'b00000000000000000000000000000000 : n2384;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2416 = n1500 ? 1'b0 : n2386;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2417 = n1500 ? n1574 : n2387;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2418 = n1500 ? fpcr : n2388;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2419 = n1500 ? fpsr : n2389;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2420 = n1500 ? n919 : n2390;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2421 = n1500 ? n1576 : n2392;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2423 = n1500 ? fsave_frame_format_latched : n2394;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2424 = n1500 ? n1577 : n2395;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2425 = n1500 ? n1578 : n2396;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2426 = n1500 ? fsave_counter : n2397;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2427 = n1500 ? frestore_frame_format : n2398;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2430 = n1500 ? n1580 : n2401;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2431 = n1500 ? converter_start : n2402;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2432 = n1500 ? converter_source_format : n2403;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2433 = n1500 ? converter_dest_format : n2404;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2434 = n1500 ? converter_data_in : n2405;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2435 = n1500 ? rom_offset : n2406;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2436 = n1500 ? rom_read_enable : n2407;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2437 = n1500 ? n1581 : movem_predecrement;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2438 = n1500 ? n1582 : movem_postincrement;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2442 = n1500 ? fp_to_int_shift : n2411;
  /* TG68K_FPU.vhd:1582:41  */
  assign n2443 = n1500 ? fp_to_int_result : n2412;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2444 = n1267 ? n1413 : n2414;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2445 = n1267 ? n1493 : n2416;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2446 = n1267 ? n1417 : n2417;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2447 = n1267 ? n1418 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2448 = n1267 ? n1419 : fp_reg_write_addr;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2449 = n1267 ? n1420 : fp_reg_write_data;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2451 = n1267 ? n1422 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2452 = n1267 ? fpcr : n2418;
  assign n2453 = n2419[27:0]; // extract
  assign n2454 = fpsr[27:0]; // extract
  /* TG68K_FPU.vhd:1499:41  */
  assign n2455 = n1267 ? n2454 : n2453;
  assign n2456 = n2419[31:28]; // extract
  /* TG68K_FPU.vhd:1499:41  */
  assign n2457 = n1267 ? n1496 : n2456;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2458 = n1267 ? n919 : n2420;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2459 = n1267 ? n1498 : n2421;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2461 = n1267 ? fsave_frame_format_latched : n2423;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2462 = n1267 ? movem_register_list : n2424;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2463 = n1267 ? movem_direction : n2425;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2464 = n1267 ? fsave_counter : n2426;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2465 = n1267 ? frestore_frame_format : n2427;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2468 = n1267 ? n1426 : n2430;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2469 = n1267 ? converter_start : n2431;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2470 = n1267 ? converter_source_format : n2432;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2471 = n1267 ? converter_dest_format : n2433;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2472 = n1267 ? converter_data_in : n2434;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2473 = n1267 ? n1427 : n2435;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2474 = n1267 ? n1429 : n2436;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2475 = n1267 ? movem_predecrement : n2437;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2476 = n1267 ? movem_postincrement : n2438;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2480 = n1267 ? fp_to_int_shift : n2442;
  /* TG68K_FPU.vhd:1499:41  */
  assign n2481 = n1267 ? fp_to_int_result : n2443;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2483 = n1215 ? 32'b00000000000000000000000000000000 : n2444;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2485 = n1215 ? 1'b0 : n2445;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2486 = n1215 ? n910 : n2446;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2487 = n1215 ? fp_reg_write_enable : n2447;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2488 = n1215 ? fp_reg_write_addr : n2448;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2489 = n1215 ? fp_reg_write_data : n2449;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2491 = n1215 ? fp_reg_access_valid : n2451;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2492 = n1215 ? fpcr : n2452;
  assign n2493 = {n2457, n2455};
  assign n2494 = n2493[27:0]; // extract
  assign n2495 = fpsr[27:0]; // extract
  /* TG68K_FPU.vhd:1457:41  */
  assign n2496 = n1215 ? n2495 : n2494;
  assign n2497 = n2493[31:28]; // extract
  /* TG68K_FPU.vhd:1457:41  */
  assign n2498 = n1215 ? n1250 : n2497;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2499 = n1215 ? n919 : n2458;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2501 = n1215 ? 4'b0101 : n2459;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2503 = n1215 ? fsave_frame_format_latched : n2461;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2504 = n1215 ? movem_register_list : n2462;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2505 = n1215 ? movem_direction : n2463;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2506 = n1215 ? fsave_counter : n2464;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2507 = n1215 ? frestore_frame_format : n2465;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2510 = n1215 ? n913 : n2468;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2511 = n1215 ? converter_start : n2469;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2512 = n1215 ? converter_source_format : n2470;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2513 = n1215 ? converter_dest_format : n2471;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2514 = n1215 ? converter_data_in : n2472;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2515 = n1215 ? rom_offset : n2473;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2516 = n1215 ? rom_read_enable : n2474;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2517 = n1215 ? movem_predecrement : n2475;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2518 = n1215 ? movem_postincrement : n2476;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2522 = n1215 ? fp_to_int_shift : n2480;
  /* TG68K_FPU.vhd:1457:41  */
  assign n2523 = n1215 ? fp_to_int_result : n2481;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2525 = n1109 ? 32'b00000000000000000000000000000000 : n2483;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2526 = n1109 ? n1200 : n2485;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2527 = n1109 ? n1202 : n2486;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2528 = n1109 ? fp_reg_write_enable : n2487;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2529 = n1109 ? fp_reg_write_addr : n2488;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2530 = n1109 ? fp_reg_write_data : n2489;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2532 = n1109 ? fp_reg_access_valid : n2491;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2533 = n1109 ? fpcr : n2492;
  assign n2534 = {n2498, n2496};
  /* TG68K_FPU.vhd:1442:41  */
  assign n2535 = n1109 ? fpsr : n2534;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2536 = n1109 ? n919 : n2499;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2537 = n1109 ? n1205 : n2501;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2539 = n1109 ? fsave_frame_format_latched : n2503;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2540 = n1109 ? movem_register_list : n2504;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2541 = n1109 ? movem_direction : n2505;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2542 = n1109 ? fsave_counter : n2506;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2543 = n1109 ? frestore_frame_format : n2507;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2546 = n1109 ? n1207 : n2510;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2547 = n1109 ? converter_start : n2511;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2548 = n1109 ? converter_source_format : n2512;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2549 = n1109 ? converter_dest_format : n2513;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2550 = n1109 ? converter_data_in : n2514;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2551 = n1109 ? rom_offset : n2515;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2552 = n1109 ? rom_read_enable : n2516;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2553 = n1109 ? movem_predecrement : n2517;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2554 = n1109 ? movem_postincrement : n2518;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2558 = n1109 ? fp_to_int_shift : n2522;
  /* TG68K_FPU.vhd:1442:41  */
  assign n2559 = n1109 ? fp_to_int_result : n2523;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2560 = n1016 ? n1107 : n2525;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2562 = n1016 ? 1'b1 : n2526;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2563 = n1016 ? n910 : n2527;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2564 = n1016 ? fp_reg_write_enable : n2528;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2565 = n1016 ? fp_reg_write_addr : n2529;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2566 = n1016 ? fp_reg_write_data : n2530;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2568 = n1016 ? fp_reg_access_valid : n2532;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2569 = n1016 ? fpcr : n2533;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2570 = n1016 ? fpsr : n2535;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2571 = n1016 ? n919 : n2536;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2573 = n1016 ? 4'b0000 : n2537;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2575 = n1016 ? fsave_frame_format_latched : n2539;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2576 = n1016 ? movem_register_list : n2540;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2577 = n1016 ? movem_direction : n2541;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2578 = n1016 ? fsave_counter : n2542;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2579 = n1016 ? frestore_frame_format : n2543;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2582 = n1016 ? n913 : n2546;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2583 = n1016 ? converter_start : n2547;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2584 = n1016 ? converter_source_format : n2548;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2585 = n1016 ? converter_dest_format : n2549;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2586 = n1016 ? converter_data_in : n2550;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2587 = n1016 ? rom_offset : n2551;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2588 = n1016 ? rom_read_enable : n2552;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2589 = n1016 ? movem_predecrement : n2553;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2590 = n1016 ? movem_postincrement : n2554;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2594 = n1016 ? fp_to_int_shift : n2558;
  /* TG68K_FPU.vhd:1431:41  */
  assign n2595 = n1016 ? fp_to_int_result : n2559;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2596 = n922 ? n1014 : n2560;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2598 = n922 ? 1'b1 : n2562;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2599 = n922 ? n910 : n2563;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2600 = n922 ? fp_reg_write_enable : n2564;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2601 = n922 ? fp_reg_write_addr : n2565;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2602 = n922 ? fp_reg_write_data : n2566;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2604 = n922 ? fp_reg_access_valid : n2568;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2605 = n922 ? fpcr : n2569;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2606 = n922 ? fpsr : n2570;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2607 = n922 ? n919 : n2571;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2609 = n922 ? 4'b0000 : n2573;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2611 = n922 ? fsave_frame_format_latched : n2575;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2612 = n922 ? movem_register_list : n2576;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2613 = n922 ? movem_direction : n2577;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2614 = n922 ? fsave_counter : n2578;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2615 = n922 ? frestore_frame_format : n2579;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2618 = n922 ? n913 : n2582;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2619 = n922 ? converter_start : n2583;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2620 = n922 ? converter_source_format : n2584;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2621 = n922 ? converter_dest_format : n2585;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2622 = n922 ? converter_data_in : n2586;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2623 = n922 ? rom_offset : n2587;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2624 = n922 ? rom_read_enable : n2588;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2625 = n922 ? movem_predecrement : n2589;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2626 = n922 ? movem_postincrement : n2590;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2630 = n922 ? fp_to_int_shift : n2594;
  /* TG68K_FPU.vhd:1417:41  */
  assign n2631 = n922 ? fp_to_int_result : n2595;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2633 = n920 ? 32'b00000000000000000000000000000000 : n2596;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2635 = n920 ? 1'b0 : n2598;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2637 = n920 ? 1'b1 : n2599;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2638 = n920 ? fp_reg_write_enable : n2600;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2639 = n920 ? fp_reg_write_addr : n2601;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2640 = n920 ? fp_reg_write_data : n2602;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2642 = n920 ? fp_reg_access_valid : n2604;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2643 = n920 ? fpcr : n2605;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2644 = n920 ? fpsr : n2606;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2645 = n920 ? n919 : n2607;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2647 = n920 ? 4'b1000 : n2609;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2649 = n920 ? fsave_frame_format_latched : n2611;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2650 = n920 ? movem_register_list : n2612;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2651 = n920 ? movem_direction : n2613;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2652 = n920 ? fsave_counter : n2614;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2653 = n920 ? frestore_frame_format : n2615;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2657 = n920 ? 8'b00010000 : n2618;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2658 = n920 ? converter_start : n2619;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2659 = n920 ? converter_source_format : n2620;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2660 = n920 ? converter_dest_format : n2621;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2661 = n920 ? converter_data_in : n2622;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2662 = n920 ? rom_offset : n2623;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2663 = n920 ? rom_read_enable : n2624;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2664 = n920 ? movem_predecrement : n2625;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2665 = n920 ? movem_postincrement : n2626;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2669 = n920 ? fp_to_int_shift : n2630;
  /* TG68K_FPU.vhd:1411:49  */
  assign n2670 = n920 ? fp_to_int_result : n2631;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2672 = decoder_unsupported ? 32'b00000000000000000000000000000000 : n2633;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2674 = decoder_unsupported ? 1'b0 : n2635;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2676 = decoder_unsupported ? 1'b1 : n2637;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2677 = decoder_unsupported ? fp_reg_write_enable : n2638;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2678 = decoder_unsupported ? fp_reg_write_addr : n2639;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2679 = decoder_unsupported ? fp_reg_write_data : n2640;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2681 = decoder_unsupported ? fp_reg_access_valid : n2642;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2682 = decoder_unsupported ? fpcr : n2643;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2683 = decoder_unsupported ? fpsr : n2644;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2684 = decoder_unsupported ? n919 : n2645;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2686 = decoder_unsupported ? 4'b1000 : n2647;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2688 = decoder_unsupported ? fsave_frame_format_latched : n2649;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2689 = decoder_unsupported ? movem_register_list : n2650;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2690 = decoder_unsupported ? movem_direction : n2651;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2691 = decoder_unsupported ? fsave_counter : n2652;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2692 = decoder_unsupported ? frestore_frame_format : n2653;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2696 = decoder_unsupported ? 8'b00001100 : n2657;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2697 = decoder_unsupported ? converter_start : n2658;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2698 = decoder_unsupported ? converter_source_format : n2659;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2699 = decoder_unsupported ? converter_dest_format : n2660;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2700 = decoder_unsupported ? converter_data_in : n2661;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2701 = decoder_unsupported ? rom_offset : n2662;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2702 = decoder_unsupported ? rom_read_enable : n2663;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2703 = decoder_unsupported ? movem_predecrement : n2664;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2704 = decoder_unsupported ? movem_postincrement : n2665;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2708 = decoder_unsupported ? fp_to_int_shift : n2669;
  /* TG68K_FPU.vhd:1406:49  */
  assign n2709 = decoder_unsupported ? fp_to_int_result : n2670;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2711 = decoder_illegal ? 32'b00000000000000000000000000000000 : n2672;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2713 = decoder_illegal ? 1'b0 : n2674;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2715 = decoder_illegal ? 1'b1 : n2676;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2716 = decoder_illegal ? fp_reg_write_enable : n2677;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2717 = decoder_illegal ? fp_reg_write_addr : n2678;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2718 = decoder_illegal ? fp_reg_write_data : n2679;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2720 = decoder_illegal ? fp_reg_access_valid : n2681;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2721 = decoder_illegal ? fpcr : n2682;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2722 = decoder_illegal ? fpsr : n2683;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2723 = decoder_illegal ? n919 : n2684;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2725 = decoder_illegal ? 4'b1000 : n2686;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2727 = decoder_illegal ? fsave_frame_format_latched : n2688;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2728 = decoder_illegal ? movem_register_list : n2689;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2729 = decoder_illegal ? movem_direction : n2690;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2730 = decoder_illegal ? fsave_counter : n2691;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2731 = decoder_illegal ? frestore_frame_format : n2692;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2735 = decoder_illegal ? 8'b00010000 : n2696;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2736 = decoder_illegal ? converter_start : n2697;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2737 = decoder_illegal ? converter_source_format : n2698;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2738 = decoder_illegal ? converter_dest_format : n2699;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2739 = decoder_illegal ? converter_data_in : n2700;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2740 = decoder_illegal ? rom_offset : n2701;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2741 = decoder_illegal ? rom_read_enable : n2702;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2742 = decoder_illegal ? movem_predecrement : n2703;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2743 = decoder_illegal ? movem_postincrement : n2704;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2747 = decoder_illegal ? fp_to_int_shift : n2708;
  /* TG68K_FPU.vhd:1401:49  */
  assign n2748 = decoder_illegal ? fp_to_int_result : n2709;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2750 = command_valid ? n2711 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2753 = command_valid ? n2713 : 1'b0;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2755 = command_valid ? n2715 : n910;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2756 = command_valid ? n2716 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2757 = command_valid ? n2717 : fp_reg_write_addr;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2758 = command_valid ? n2718 : fp_reg_write_data;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2760 = command_valid ? n2720 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2761 = command_valid ? n2721 : fpcr;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2762 = command_valid ? n2722 : fpsr;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2763 = command_valid ? n2723 : fpiar;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2764 = command_valid ? opcode : operation_word_cir;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2765 = command_valid ? cpu_address_in : command_address_cir;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2766 = command_valid ? n2725 : n912;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2768 = command_valid ? n2727 : fsave_frame_format_latched;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2769 = command_valid ? n2728 : movem_register_list;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2770 = command_valid ? n2729 : movem_direction;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2771 = command_valid ? n2730 : fsave_counter;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2772 = command_valid ? n2731 : frestore_frame_format;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2775 = command_valid ? n2735 : n913;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2776 = command_valid ? n2736 : converter_start;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2777 = command_valid ? n2737 : converter_source_format;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2778 = command_valid ? n2738 : converter_dest_format;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2779 = command_valid ? n2739 : converter_data_in;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2780 = command_valid ? n2740 : rom_offset;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2781 = command_valid ? n2741 : rom_read_enable;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2782 = command_valid ? n2742 : movem_predecrement;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2783 = command_valid ? n2743 : movem_postincrement;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2787 = command_valid ? n2747 : fp_to_int_shift;
  /* TG68K_FPU.vhd:1384:49  */
  assign n2788 = command_valid ? n2748 : fp_to_int_result;
  /* TG68K_FPU.vhd:1306:41  */
  assign n2790 = fpu_state == 4'b0001;
  /* TG68K_FPU.vhd:2095:67  */
  assign n2792 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:2095:94  */
  assign n2794 = fpu_operation == 7'b0111000;
  /* TG68K_FPU.vhd:2095:77  */
  assign n2795 = n2792 | n2794;
  /* TG68K_FPU.vhd:2095:105  */
  assign n2796 = cir_write & n2795;
  /* TG68K_FPU.vhd:2096:84  */
  assign n2798 = cir_address == 5'b00101;
  /* TG68K_FPU.vhd:2096:68  */
  assign n2799 = n2798 & n2796;
  /* TG68K_FPU.vhd:2102:87  */
  assign n2800 = cir_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2102:100  */
  assign n2802 = n2800 == 8'b00000000;
  /* TG68K_FPU.vhd:2105:90  */
  assign n2803 = cir_data_in[7]; // extract
  /* TG68K_FPU.vhd:2105:94  */
  assign n2804 = ~n2803;
  /* TG68K_FPU.vhd:2107:95  */
  assign n2805 = cir_data_in[6]; // extract
  /* TG68K_FPU.vhd:2109:116  */
  assign n2806 = cir_data_in[6:0]; // extract
  /* TG68K_FPU.vhd:2108:159  */
  assign n2808 = {17'b01000000000001011, n2806};
  /* TG68K_FPU.vhd:2109:129  */
  assign n2810 = {n2808, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2110:98  */
  assign n2811 = cir_data_in[5]; // extract
  /* TG68K_FPU.vhd:2112:116  */
  assign n2812 = cir_data_in[5:0]; // extract
  /* TG68K_FPU.vhd:2111:159  */
  assign n2814 = {17'b01000000000001001, n2812};
  /* TG68K_FPU.vhd:2112:129  */
  assign n2816 = {n2814, 1'b0};
  /* TG68K_FPU.vhd:2112:135  */
  assign n2818 = {n2816, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2113:98  */
  assign n2819 = cir_data_in[4]; // extract
  /* TG68K_FPU.vhd:2115:116  */
  assign n2820 = cir_data_in[4:0]; // extract
  /* TG68K_FPU.vhd:2114:159  */
  assign n2822 = {17'b01000000000000111, n2820};
  /* TG68K_FPU.vhd:2115:129  */
  assign n2824 = {n2822, 2'b00};
  /* TG68K_FPU.vhd:2115:136  */
  assign n2826 = {n2824, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2116:98  */
  assign n2827 = cir_data_in[3]; // extract
  /* TG68K_FPU.vhd:2118:116  */
  assign n2828 = cir_data_in[3:0]; // extract
  /* TG68K_FPU.vhd:2117:159  */
  assign n2830 = {17'b01000000000000101, n2828};
  /* TG68K_FPU.vhd:2118:129  */
  assign n2832 = {n2830, 3'b000};
  /* TG68K_FPU.vhd:2118:137  */
  assign n2834 = {n2832, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2119:98  */
  assign n2835 = cir_data_in[2]; // extract
  /* TG68K_FPU.vhd:2121:116  */
  assign n2836 = cir_data_in[2:0]; // extract
  /* TG68K_FPU.vhd:2120:159  */
  assign n2838 = {17'b01000000000000011, n2836};
  /* TG68K_FPU.vhd:2121:129  */
  assign n2840 = {n2838, 4'b0000};
  /* TG68K_FPU.vhd:2121:138  */
  assign n2842 = {n2840, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2122:98  */
  assign n2843 = cir_data_in[1]; // extract
  /* TG68K_FPU.vhd:2124:116  */
  assign n2844 = cir_data_in[1:0]; // extract
  /* TG68K_FPU.vhd:2123:159  */
  assign n2846 = {17'b01000000000000001, n2844};
  /* TG68K_FPU.vhd:2124:129  */
  assign n2848 = {n2846, 5'b00000};
  /* TG68K_FPU.vhd:2124:139  */
  assign n2850 = {n2848, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2127:116  */
  assign n2851 = cir_data_in[0]; // extract
  /* TG68K_FPU.vhd:2126:159  */
  assign n2853 = {17'b00111111111111111, n2851};
  /* TG68K_FPU.vhd:2127:129  */
  assign n2855 = {n2853, 6'b000000};
  /* TG68K_FPU.vhd:2127:140  */
  assign n2857 = {n2855, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2122:81  */
  assign n2858 = n2843 ? n2850 : n2857;
  /* TG68K_FPU.vhd:2119:81  */
  assign n2859 = n2835 ? n2842 : n2858;
  /* TG68K_FPU.vhd:2116:81  */
  assign n2860 = n2827 ? n2834 : n2859;
  /* TG68K_FPU.vhd:2113:81  */
  assign n2861 = n2819 ? n2826 : n2860;
  /* TG68K_FPU.vhd:2110:81  */
  assign n2862 = n2811 ? n2818 : n2861;
  /* TG68K_FPU.vhd:2107:81  */
  assign n2863 = n2805 ? n2810 : n2862;
  /* TG68K_FPU.vhd:2131:95  */
  assign n2864 = cir_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2131:108  */
  assign n2866 = n2864 == 8'b10000000;
  /* TG68K_FPU.vhd:2139:147  */
  assign n2867 = cir_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2139:132  */
  assign n2868 = ~n2867;
  /* TG68K_FPU.vhd:2139:161  */
  assign n2870 = n2868 + 8'b00000001;
  /* TG68K_FPU.vhd:2138:163  */
  assign n2872 = {17'b11000000000001101, n2870};
  /* TG68K_FPU.vhd:2139:167  */
  assign n2874 = {n2872, 55'b0000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2131:81  */
  assign n2876 = n2866 ? 80'b11000000000001101100000000000000000000000000000000000000000000000000000000000000 : n2874;
  /* TG68K_FPU.vhd:2105:73  */
  assign n2877 = n2804 ? n2863 : n2876;
  /* TG68K_FPU.vhd:2102:73  */
  assign n2879 = n2802 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n2877;
  /* TG68K_FPU.vhd:2100:65  */
  assign n2881 = decoder_source_format == 3'b110;
  /* TG68K_FPU.vhd:2145:101  */
  assign n2883 = cir_data_in == 16'b0000000000000000;
  /* TG68K_FPU.vhd:2147:90  */
  assign n2884 = cir_data_in[15]; // extract
  /* TG68K_FPU.vhd:2147:95  */
  assign n2885 = ~n2884;
  /* TG68K_FPU.vhd:2149:122  */
  assign n2887 = {16'b0100000000001110, cir_data_in};
  /* TG68K_FPU.vhd:2149:149  */
  assign n2889 = {n2887, 48'b000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2152:126  */
  assign n2890 = ~cir_data_in;
  /* TG68K_FPU.vhd:2152:156  */
  assign n2892 = n2890 + 16'b0000000000000001;
  /* TG68K_FPU.vhd:2152:122  */
  assign n2894 = {16'b1100000000001110, n2892};
  /* TG68K_FPU.vhd:2152:161  */
  assign n2896 = {n2894, 48'b000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2147:73  */
  assign n2897 = n2885 ? n2889 : n2896;
  /* TG68K_FPU.vhd:2145:73  */
  assign n2899 = n2883 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n2897;
  /* TG68K_FPU.vhd:2143:65  */
  assign n2901 = decoder_source_format == 3'b100;
  /* TG68K_FPU.vhd:2158:120  */
  assign n2903 = {17'b00111111100000001, cir_data_in};
  /* TG68K_FPU.vhd:2158:147  */
  assign n2905 = {n2903, 47'b00000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2155:65  */
  assign n2907 = decoder_source_format == 3'b000;
  assign n2908 = {n2907, n2901, n2881};
  /* TG68K_FPU.vhd:2099:57  */
  always @*
    case (n2908)
      3'b100: n2910 = n2905;
      3'b010: n2910 = n2899;
      3'b001: n2910 = n2879;
      default: n2910 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:2167:70  */
  assign n2912 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:2167:97  */
  assign n2914 = fpu_operation == 7'b0111000;
  /* TG68K_FPU.vhd:2167:80  */
  assign n2915 = n2912 | n2914;
  /* TG68K_FPU.vhd:2174:52  */
  assign n2916 = {28'b0, source_reg};  //  uext
  /* TG68K_FPU.vhd:2174:85  */
  assign n2917 = {1'b0, n2916};  //  uext
  /* TG68K_FPU.vhd:2174:85  */
  assign n2919 = $signed(n2917) > $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:2180:87  */
  assign n2922 = 3'b111 - source_reg;
  /* TG68K_FPU.vhd:2174:49  */
  assign n2926 = n2919 ? 1'b1 : fpu_exception_i;
  /* TG68K_FPU.vhd:2174:49  */
  assign n2928 = n2919 ? 4'b1000 : fpu_state;
  /* TG68K_FPU.vhd:2174:49  */
  assign n2930 = n2919 ? 8'b00001100 : exception_code_internal;
  /* TG68K_FPU.vhd:2174:49  */
  assign n2931 = n2919 ? alu_operand_a : n6960;
  /* TG68K_FPU.vhd:2182:60  */
  assign n2933 = ea_mode == 3'b000;
  /* TG68K_FPU.vhd:2190:87  */
  assign n2934 = cpu_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2190:100  */
  assign n2936 = n2934 == 8'b00000000;
  /* TG68K_FPU.vhd:2193:90  */
  assign n2937 = cpu_data_in[7]; // extract
  /* TG68K_FPU.vhd:2193:94  */
  assign n2938 = ~n2937;
  /* TG68K_FPU.vhd:2196:95  */
  assign n2939 = cpu_data_in[6]; // extract
  /* TG68K_FPU.vhd:2200:116  */
  assign n2940 = cpu_data_in[6:0]; // extract
  /* TG68K_FPU.vhd:2199:159  */
  assign n2942 = {17'b01000000000001011, n2940};
  /* TG68K_FPU.vhd:2200:129  */
  assign n2944 = {n2942, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2201:98  */
  assign n2945 = cpu_data_in[5]; // extract
  /* TG68K_FPU.vhd:2205:116  */
  assign n2946 = cpu_data_in[5:0]; // extract
  /* TG68K_FPU.vhd:2204:159  */
  assign n2948 = {17'b01000000000001001, n2946};
  /* TG68K_FPU.vhd:2205:129  */
  assign n2950 = {n2948, 1'b0};
  /* TG68K_FPU.vhd:2205:135  */
  assign n2952 = {n2950, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2206:98  */
  assign n2953 = cpu_data_in[4]; // extract
  /* TG68K_FPU.vhd:2210:116  */
  assign n2954 = cpu_data_in[4:0]; // extract
  /* TG68K_FPU.vhd:2209:159  */
  assign n2956 = {17'b01000000000000111, n2954};
  /* TG68K_FPU.vhd:2210:129  */
  assign n2958 = {n2956, 2'b00};
  /* TG68K_FPU.vhd:2210:136  */
  assign n2960 = {n2958, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2211:98  */
  assign n2961 = cpu_data_in[3]; // extract
  /* TG68K_FPU.vhd:2215:116  */
  assign n2962 = cpu_data_in[3:0]; // extract
  /* TG68K_FPU.vhd:2214:159  */
  assign n2964 = {17'b01000000000000101, n2962};
  /* TG68K_FPU.vhd:2215:129  */
  assign n2966 = {n2964, 3'b000};
  /* TG68K_FPU.vhd:2215:137  */
  assign n2968 = {n2966, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2216:98  */
  assign n2969 = cpu_data_in[2]; // extract
  /* TG68K_FPU.vhd:2220:116  */
  assign n2970 = cpu_data_in[2:0]; // extract
  /* TG68K_FPU.vhd:2219:159  */
  assign n2972 = {17'b01000000000000011, n2970};
  /* TG68K_FPU.vhd:2220:129  */
  assign n2974 = {n2972, 4'b0000};
  /* TG68K_FPU.vhd:2220:138  */
  assign n2976 = {n2974, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2221:98  */
  assign n2977 = cpu_data_in[1]; // extract
  /* TG68K_FPU.vhd:2225:116  */
  assign n2978 = cpu_data_in[1:0]; // extract
  /* TG68K_FPU.vhd:2224:159  */
  assign n2980 = {17'b01000000000000001, n2978};
  /* TG68K_FPU.vhd:2225:129  */
  assign n2982 = {n2980, 5'b00000};
  /* TG68K_FPU.vhd:2225:139  */
  assign n2984 = {n2982, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2230:116  */
  assign n2985 = cpu_data_in[0]; // extract
  /* TG68K_FPU.vhd:2229:159  */
  assign n2987 = {17'b00111111111111111, n2985};
  /* TG68K_FPU.vhd:2230:129  */
  assign n2989 = {n2987, 6'b000000};
  /* TG68K_FPU.vhd:2230:140  */
  assign n2991 = {n2989, 56'b00000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2221:81  */
  assign n2992 = n2977 ? n2984 : n2991;
  /* TG68K_FPU.vhd:2216:81  */
  assign n2993 = n2969 ? n2976 : n2992;
  /* TG68K_FPU.vhd:2211:81  */
  assign n2994 = n2961 ? n2968 : n2993;
  /* TG68K_FPU.vhd:2206:81  */
  assign n2995 = n2953 ? n2960 : n2994;
  /* TG68K_FPU.vhd:2201:81  */
  assign n2996 = n2945 ? n2952 : n2995;
  /* TG68K_FPU.vhd:2196:81  */
  assign n2997 = n2939 ? n2944 : n2996;
  /* TG68K_FPU.vhd:2234:95  */
  assign n2998 = cpu_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2234:108  */
  assign n3000 = n2998 == 8'b10000000;
  /* TG68K_FPU.vhd:2242:147  */
  assign n3001 = cpu_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2242:132  */
  assign n3002 = ~n3001;
  /* TG68K_FPU.vhd:2242:161  */
  assign n3004 = n3002 + 8'b00000001;
  /* TG68K_FPU.vhd:2241:163  */
  assign n3006 = {17'b11000000000001101, n3004};
  /* TG68K_FPU.vhd:2242:167  */
  assign n3008 = {n3006, 55'b0000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2234:81  */
  assign n3010 = n3000 ? 80'b11000000000001101100000000000000000000000000000000000000000000000000000000000000 : n3008;
  /* TG68K_FPU.vhd:2193:73  */
  assign n3011 = n2938 ? n2997 : n3010;
  /* TG68K_FPU.vhd:2190:73  */
  assign n3013 = n2936 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3011;
  /* TG68K_FPU.vhd:2186:65  */
  assign n3015 = data_format == 3'b110;
  /* TG68K_FPU.vhd:2247:87  */
  assign n3016 = cpu_data_in[15:0]; // extract
  /* TG68K_FPU.vhd:2247:101  */
  assign n3018 = n3016 == 16'b0000000000000000;
  /* TG68K_FPU.vhd:2250:90  */
  assign n3019 = cpu_data_in[15]; // extract
  /* TG68K_FPU.vhd:2250:95  */
  assign n3020 = ~n3019;
  /* TG68K_FPU.vhd:2252:135  */
  assign n3021 = cpu_data_in[15:0]; // extract
  /* TG68K_FPU.vhd:2252:122  */
  assign n3023 = {16'b0100000000001110, n3021};
  /* TG68K_FPU.vhd:2252:149  */
  assign n3025 = {n3023, 48'b000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2255:141  */
  assign n3026 = cpu_data_in[15:0]; // extract
  /* TG68K_FPU.vhd:2255:126  */
  assign n3027 = ~n3026;
  /* TG68K_FPU.vhd:2255:156  */
  assign n3029 = n3027 + 16'b0000000000000001;
  /* TG68K_FPU.vhd:2255:122  */
  assign n3031 = {16'b1100000000001110, n3029};
  /* TG68K_FPU.vhd:2255:161  */
  assign n3033 = {n3031, 48'b000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2250:73  */
  assign n3034 = n3020 ? n3025 : n3033;
  /* TG68K_FPU.vhd:2247:73  */
  assign n3036 = n3018 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3034;
  /* TG68K_FPU.vhd:2245:65  */
  assign n3038 = data_format == 3'b100;
  /* TG68K_FPU.vhd:2259:88  */
  assign n3040 = cpu_data_in == 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:2262:90  */
  assign n3041 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2262:95  */
  assign n3042 = ~n3041;
  /* TG68K_FPU.vhd:2264:122  */
  assign n3044 = {16'b0100000000011110, cpu_data_in};
  /* TG68K_FPU.vhd:2264:136  */
  assign n3046 = {n3044, 32'b00000000000000000000000000000000};
  /* TG68K_FPU.vhd:2267:126  */
  assign n3047 = ~cpu_data_in;
  /* TG68K_FPU.vhd:2267:143  */
  assign n3049 = n3047 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:2267:122  */
  assign n3051 = {16'b1100000000011110, n3049};
  /* TG68K_FPU.vhd:2267:148  */
  assign n3053 = {n3051, 32'b00000000000000000000000000000000};
  /* TG68K_FPU.vhd:2262:73  */
  assign n3054 = n3042 ? n3046 : n3053;
  /* TG68K_FPU.vhd:2259:73  */
  assign n3056 = n3040 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3054;
  /* TG68K_FPU.vhd:2257:65  */
  assign n3058 = data_format == 3'b000;
  assign n3059 = {n3058, n3038, n3015};
  /* TG68K_FPU.vhd:2185:57  */
  always @*
    case (n3059)
      3'b100: n3061 = n3056;
      3'b010: n3061 = n3036;
      3'b001: n3061 = n3013;
      default: n3061 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:2276:65  */
  assign n3063 = ea_mode == 3'b000;
  /* TG68K_FPU.vhd:2278:65  */
  assign n3065 = ea_mode == 3'b001;
  /* TG68K_FPU.vhd:2280:65  */
  assign n3067 = ea_mode == 3'b010;
  /* TG68K_FPU.vhd:2286:65  */
  assign n3069 = ea_mode == 3'b011;
  /* TG68K_FPU.vhd:2292:65  */
  assign n3071 = ea_mode == 3'b100;
  /* TG68K_FPU.vhd:2299:65  */
  assign n3073 = ea_mode == 3'b101;
  /* TG68K_FPU.vhd:2305:65  */
  assign n3075 = ea_mode == 3'b110;
  /* TG68K_FPU.vhd:2313:81  */
  assign n3077 = ea_register == 3'b000;
  /* TG68K_FPU.vhd:2319:81  */
  assign n3079 = ea_register == 3'b001;
  /* TG68K_FPU.vhd:2325:81  */
  assign n3081 = ea_register == 3'b010;
  /* TG68K_FPU.vhd:2331:81  */
  assign n3083 = ea_register == 3'b011;
  /* TG68K_FPU.vhd:2342:119  */
  assign n3084 = cpu_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2342:132  */
  assign n3086 = n3084 == 8'b00000000;
  /* TG68K_FPU.vhd:2344:122  */
  assign n3087 = cpu_data_in[7]; // extract
  /* TG68K_FPU.vhd:2344:126  */
  assign n3088 = ~n3087;
  /* TG68K_FPU.vhd:2346:157  */
  assign n3089 = cpu_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2346:144  */
  assign n3091 = {17'b00100000000000110, n3089};
  /* TG68K_FPU.vhd:2346:170  */
  assign n3093 = {n3091, 52'b0000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2346:189  */
  assign n3095 = {n3093, 3'b000};
  /* TG68K_FPU.vhd:2349:162  */
  assign n3096 = cpu_data_in[7:0]; // extract
  /* TG68K_FPU.vhd:2349:147  */
  assign n3097 = ~n3096;
  /* TG68K_FPU.vhd:2349:144  */
  assign n3099 = {17'b10100000000000110, n3097};
  /* TG68K_FPU.vhd:2349:176  */
  assign n3101 = n3099 + 25'b0000000000000000000000001;
  /* TG68K_FPU.vhd:2349:180  */
  assign n3103 = {n3101, 52'b0000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2349:199  */
  assign n3105 = {n3103, 3'b000};
  /* TG68K_FPU.vhd:2344:105  */
  assign n3106 = n3088 ? n3095 : n3105;
  /* TG68K_FPU.vhd:2342:105  */
  assign n3108 = n3086 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3106;
  /* TG68K_FPU.vhd:2340:97  */
  assign n3110 = data_format == 3'b110;
  /* TG68K_FPU.vhd:2353:119  */
  assign n3111 = cpu_data_in[15:0]; // extract
  /* TG68K_FPU.vhd:2353:133  */
  assign n3113 = n3111 == 16'b0000000000000000;
  /* TG68K_FPU.vhd:2355:122  */
  assign n3114 = cpu_data_in[15]; // extract
  /* TG68K_FPU.vhd:2355:127  */
  assign n3115 = ~n3114;
  /* TG68K_FPU.vhd:2357:157  */
  assign n3116 = cpu_data_in[15:0]; // extract
  /* TG68K_FPU.vhd:2357:144  */
  assign n3118 = {17'b00100000000001110, n3116};
  /* TG68K_FPU.vhd:2357:171  */
  assign n3120 = {n3118, 44'b00000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2357:188  */
  assign n3122 = {n3120, 3'b111};
  /* TG68K_FPU.vhd:2360:162  */
  assign n3123 = cpu_data_in[15:0]; // extract
  /* TG68K_FPU.vhd:2360:147  */
  assign n3124 = ~n3123;
  /* TG68K_FPU.vhd:2360:144  */
  assign n3126 = {17'b10100000000001110, n3124};
  /* TG68K_FPU.vhd:2360:177  */
  assign n3128 = n3126 + 33'b000000000000000000000000000000001;
  /* TG68K_FPU.vhd:2360:181  */
  assign n3130 = {n3128, 44'b00000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2360:198  */
  assign n3132 = {n3130, 3'b111};
  /* TG68K_FPU.vhd:2355:105  */
  assign n3133 = n3115 ? n3122 : n3132;
  /* TG68K_FPU.vhd:2353:105  */
  assign n3135 = n3113 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3133;
  /* TG68K_FPU.vhd:2351:97  */
  assign n3137 = data_format == 3'b100;
  /* TG68K_FPU.vhd:2364:120  */
  assign n3139 = cpu_data_in == 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:2366:122  */
  assign n3140 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2366:127  */
  assign n3141 = ~n3140;
  /* TG68K_FPU.vhd:2368:144  */
  assign n3143 = {17'b00100000000011110, cpu_data_in};
  /* TG68K_FPU.vhd:2368:158  */
  assign n3145 = {n3143, 28'b0000000000000000000000000000};
  /* TG68K_FPU.vhd:2368:171  */
  assign n3147 = {n3145, 3'b000};
  /* TG68K_FPU.vhd:2371:147  */
  assign n3148 = ~cpu_data_in;
  /* TG68K_FPU.vhd:2371:144  */
  assign n3150 = {17'b10100000000011110, n3148};
  /* TG68K_FPU.vhd:2371:164  */
  assign n3152 = n3150 + 49'b0000000000000000000000000000000000000000000000001;
  /* TG68K_FPU.vhd:2371:168  */
  assign n3154 = {n3152, 28'b0000000000000000000000000000};
  /* TG68K_FPU.vhd:2371:181  */
  assign n3156 = {n3154, 3'b000};
  /* TG68K_FPU.vhd:2366:105  */
  assign n3157 = n3141 ? n3147 : n3156;
  /* TG68K_FPU.vhd:2364:105  */
  assign n3159 = n3139 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3157;
  /* TG68K_FPU.vhd:2362:97  */
  assign n3161 = data_format == 3'b000;
  /* TG68K_FPU.vhd:2377:119  */
  assign n3162 = cpu_data_in[30:23]; // extract
  /* TG68K_FPU.vhd:2377:134  */
  assign n3164 = n3162 == 8'b00000000;
  /* TG68K_FPU.vhd:2379:127  */
  assign n3165 = cpu_data_in[22:0]; // extract
  /* TG68K_FPU.vhd:2379:141  */
  assign n3167 = n3165 == 23'b00000000000000000000000;
  /* TG68K_FPU.vhd:2381:149  */
  assign n3168 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2381:154  */
  assign n3170 = {n3168, 15'b000000000000000};
  /* TG68K_FPU.vhd:2381:174  */
  assign n3172 = {n3170, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2386:149  */
  assign n3173 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2386:154  */
  assign n3175 = {n3173, 16'b0011111110000001};
  /* TG68K_FPU.vhd:2386:164  */
  assign n3177 = {n3175, 1'b0};
  /* TG68K_FPU.vhd:2386:183  */
  assign n3178 = cpu_data_in[22:0]; // extract
  /* TG68K_FPU.vhd:2386:170  */
  assign n3179 = {n3177, n3178};
  /* TG68K_FPU.vhd:2386:197  */
  assign n3181 = {n3179, 36'b000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2386:212  */
  assign n3183 = {n3181, 3'b000};
  /* TG68K_FPU.vhd:2379:113  */
  assign n3184 = n3167 ? n3172 : n3183;
  /* TG68K_FPU.vhd:2388:122  */
  assign n3185 = cpu_data_in[30:23]; // extract
  /* TG68K_FPU.vhd:2388:137  */
  assign n3187 = n3185 == 8'b11111111;
  /* TG68K_FPU.vhd:2390:127  */
  assign n3188 = cpu_data_in[22:0]; // extract
  /* TG68K_FPU.vhd:2390:141  */
  assign n3190 = n3188 == 23'b00000000000000000000000;
  /* TG68K_FPU.vhd:2392:149  */
  assign n3191 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2392:154  */
  assign n3193 = {n3191, 15'b111111111111111};
  /* TG68K_FPU.vhd:2392:174  */
  assign n3195 = {n3193, 64'b1000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2395:149  */
  assign n3196 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2395:154  */
  assign n3198 = {n3196, 15'b111111111111111};
  /* TG68K_FPU.vhd:2395:174  */
  assign n3200 = {n3198, 1'b1};
  /* TG68K_FPU.vhd:2395:193  */
  assign n3201 = cpu_data_in[22:0]; // extract
  /* TG68K_FPU.vhd:2395:180  */
  assign n3202 = {n3200, n3201};
  /* TG68K_FPU.vhd:2395:207  */
  assign n3204 = {n3202, 40'b0000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2390:113  */
  assign n3205 = n3190 ? n3195 : n3204;
  /* TG68K_FPU.vhd:2400:141  */
  assign n3206 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2400:146  */
  assign n3208 = {n3206, 15'b011111110000000};
  /* TG68K_FPU.vhd:2400:166  */
  assign n3210 = {n3208, 1'b1};
  /* TG68K_FPU.vhd:2400:185  */
  assign n3211 = cpu_data_in[22:0]; // extract
  /* TG68K_FPU.vhd:2400:172  */
  assign n3212 = {n3210, n3211};
  /* TG68K_FPU.vhd:2400:199  */
  assign n3214 = {n3212, 40'b0000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2388:105  */
  assign n3215 = n3187 ? n3205 : n3214;
  /* TG68K_FPU.vhd:2377:105  */
  assign n3216 = n3164 ? n3184 : n3215;
  /* TG68K_FPU.vhd:2373:97  */
  assign n3218 = data_format == 3'b001;
  /* TG68K_FPU.vhd:2405:119  */
  assign n3219 = cpu_data_in[30:20]; // extract
  /* TG68K_FPU.vhd:2405:134  */
  assign n3221 = n3219 == 11'b00000000000;
  /* TG68K_FPU.vhd:2407:141  */
  assign n3222 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2407:146  */
  assign n3224 = {n3222, 15'b000000000000000};
  /* TG68K_FPU.vhd:2407:166  */
  assign n3226 = {n3224, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2408:122  */
  assign n3227 = cpu_data_in[30:20]; // extract
  /* TG68K_FPU.vhd:2408:137  */
  assign n3229 = n3227 == 11'b11111111111;
  /* TG68K_FPU.vhd:2410:141  */
  assign n3230 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2410:146  */
  assign n3232 = {n3230, 15'b111111111111111};
  /* TG68K_FPU.vhd:2410:179  */
  assign n3233 = cpu_data_in[19:0]; // extract
  /* TG68K_FPU.vhd:2410:166  */
  assign n3234 = {n3232, n3233};
  /* TG68K_FPU.vhd:2410:193  */
  assign n3236 = {n3234, 44'b00000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2414:141  */
  assign n3237 = cpu_data_in[31]; // extract
  /* TG68K_FPU.vhd:2414:146  */
  assign n3239 = {n3237, 15'b011110000000000};
  /* TG68K_FPU.vhd:2414:166  */
  assign n3241 = {n3239, 1'b1};
  /* TG68K_FPU.vhd:2414:185  */
  assign n3242 = cpu_data_in[19:0]; // extract
  /* TG68K_FPU.vhd:2414:172  */
  assign n3243 = {n3241, n3242};
  /* TG68K_FPU.vhd:2414:199  */
  assign n3245 = {n3243, 43'b0000000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2408:105  */
  assign n3246 = n3229 ? n3236 : n3245;
  /* TG68K_FPU.vhd:2405:105  */
  assign n3247 = n3221 ? n3226 : n3246;
  /* TG68K_FPU.vhd:2402:97  */
  assign n3249 = data_format == 3'b101;
  assign n3250 = {n3249, n3218, n3161, n3137, n3110};
  /* TG68K_FPU.vhd:2339:89  */
  always @*
    case (n3250)
      5'b10000: n3252 = n3247;
      5'b01000: n3252 = n3216;
      5'b00100: n3252 = n3159;
      5'b00010: n3252 = n3135;
      5'b00001: n3252 = n3108;
      default: n3252 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:2337:81  */
  assign n3255 = ea_register == 3'b100;
  /* TG68K_FPU.vhd:2431:81  */
  assign n3257 = ea_register == 3'b101;
  /* TG68K_FPU.vhd:2437:81  */
  assign n3259 = ea_register == 3'b110;
  /* TG68K_FPU.vhd:2443:81  */
  assign n3261 = ea_register == 3'b111;
  assign n3262 = {n3261, n3259, n3257, n3255, n3083, n3081, n3079, n3077};
  /* TG68K_FPU.vhd:2312:73  */
  always @*
    case (n3262)
      8'b10000000: n3272 = 4'b0011;
      8'b01000000: n3272 = 4'b0011;
      8'b00100000: n3272 = 4'b0011;
      8'b00010000: n3272 = 4'b0101;
      8'b00001000: n3272 = 4'b0011;
      8'b00000100: n3272 = 4'b0011;
      8'b00000010: n3272 = 4'b0011;
      8'b00000001: n3272 = 4'b0011;
      default: n3272 = 4'b0101;
    endcase
  /* TG68K_FPU.vhd:2312:73  */
  always @*
    case (n3262)
      8'b10000000: n3276 = 1'b0;
      8'b01000000: n3276 = 1'b0;
      8'b00100000: n3276 = 1'b0;
      8'b00010000: n3276 = 1'b1;
      8'b00001000: n3276 = 1'b0;
      8'b00000100: n3276 = 1'b0;
      8'b00000010: n3276 = 1'b0;
      8'b00000001: n3276 = 1'b0;
      default: n3276 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:2312:73  */
  always @*
    case (n3262)
      8'b10000000: n3277 = alu_operation_code;
      8'b01000000: n3277 = alu_operation_code;
      8'b00100000: n3277 = alu_operation_code;
      8'b00010000: n3277 = fpu_operation;
      8'b00001000: n3277 = alu_operation_code;
      8'b00000100: n3277 = alu_operation_code;
      8'b00000010: n3277 = alu_operation_code;
      8'b00000001: n3277 = alu_operation_code;
      default: n3277 = fpu_operation;
    endcase
  /* TG68K_FPU.vhd:2312:73  */
  always @*
    case (n3262)
      8'b10000000: n3279 = alu_operand_b;
      8'b01000000: n3279 = alu_operand_b;
      8'b00100000: n3279 = alu_operand_b;
      8'b00010000: n3279 = n3252;
      8'b00001000: n3279 = alu_operand_b;
      8'b00000100: n3279 = alu_operand_b;
      8'b00000010: n3279 = alu_operand_b;
      8'b00000001: n3279 = alu_operand_b;
      default: n3279 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:2311:65  */
  assign n3281 = ea_mode == 3'b111;
  assign n3282 = {n3281, n3075, n3073, n3071, n3069, n3067, n3065, n3063};
  /* TG68K_FPU.vhd:2275:57  */
  always @*
    case (n3282)
      8'b10000000: n3289 = n3272;
      8'b01000000: n3289 = 4'b0011;
      8'b00100000: n3289 = 4'b0011;
      8'b00010000: n3289 = 4'b0011;
      8'b00001000: n3289 = 4'b0011;
      8'b00000100: n3289 = 4'b0011;
      8'b00000010: n3289 = n2928;
      8'b00000001: n3289 = n2928;
      default: n3289 = 4'b0101;
    endcase
  /* TG68K_FPU.vhd:2275:57  */
  always @*
    case (n3282)
      8'b10000000: n3292 = n3276;
      8'b01000000: n3292 = 1'b0;
      8'b00100000: n3292 = 1'b0;
      8'b00010000: n3292 = 1'b0;
      8'b00001000: n3292 = 1'b0;
      8'b00000100: n3292 = 1'b0;
      8'b00000010: n3292 = 1'b0;
      8'b00000001: n3292 = 1'b0;
      default: n3292 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:2275:57  */
  always @*
    case (n3282)
      8'b10000000: n3293 = n3277;
      8'b01000000: n3293 = alu_operation_code;
      8'b00100000: n3293 = alu_operation_code;
      8'b00010000: n3293 = alu_operation_code;
      8'b00001000: n3293 = alu_operation_code;
      8'b00000100: n3293 = alu_operation_code;
      8'b00000010: n3293 = alu_operation_code;
      8'b00000001: n3293 = alu_operation_code;
      default: n3293 = fpu_operation;
    endcase
  /* TG68K_FPU.vhd:2275:57  */
  always @*
    case (n3282)
      8'b10000000: n3297 = n3279;
      8'b01000000: n3297 = alu_operand_b;
      8'b00100000: n3297 = alu_operand_b;
      8'b00010000: n3297 = alu_operand_b;
      8'b00001000: n3297 = alu_operand_b;
      8'b00000100: n3297 = alu_operand_b;
      8'b00000010: n3297 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
      8'b00000001: n3297 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
      default: n3297 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:2182:49  */
  assign n3298 = n2933 ? n2928 : n3289;
  /* TG68K_FPU.vhd:2182:49  */
  assign n3300 = n2933 ? 1'b0 : n3292;
  /* TG68K_FPU.vhd:2182:49  */
  assign n3301 = n2933 ? alu_operation_code : n3293;
  /* TG68K_FPU.vhd:2182:49  */
  assign n3302 = n2933 ? n3061 : n3297;
  /* TG68K_FPU.vhd:2466:66  */
  assign n3304 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:2466:88  */
  assign n3306 = ea_mode == 3'b111;
  /* TG68K_FPU.vhd:2466:76  */
  assign n3307 = n3306 & n3304;
  /* TG68K_FPU.vhd:2466:112  */
  assign n3309 = ea_register == 3'b010;
  /* TG68K_FPU.vhd:2466:96  */
  assign n3310 = n3309 & n3307;
  /* TG68K_FPU.vhd:550:33  */
  assign n3317 = alu_operand_a[79]; // extract
  /* TG68K_FPU.vhd:551:37  */
  assign n3319 = alu_operand_a[78:64]; // extract
  /* TG68K_FPU.vhd:552:37  */
  assign n3321 = alu_operand_a[63:0]; // extract
  /* TG68K_FPU.vhd:558:29  */
  assign n3325 = n3319 == 15'b111111111111111;
  /* TG68K_FPU.vhd:560:36  */
  assign n3326 = alu_operand_a[63]; // extract
  /* TG68K_FPU.vhd:560:41  */
  assign n3327 = ~n3326;
  /* TG68K_FPU.vhd:560:58  */
  assign n3328 = alu_operand_a[62:0]; // extract
  /* TG68K_FPU.vhd:560:72  */
  assign n3330 = n3328 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:560:47  */
  assign n3331 = n3327 | n3330;
  assign n3334 = n3323[0]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3335 = n3331 ? 1'b1 : n3334;
  assign n3336 = n3323[1]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3337 = n3331 ? n3336 : 1'b1;
  assign n3338 = n3323[3]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3339 = n3331 ? n3338 : n3317;
  /* TG68K_FPU.vhd:568:32  */
  assign n3341 = n3319 == 15'b000000000000000;
  /* TG68K_FPU.vhd:568:68  */
  assign n3343 = n3321 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:568:55  */
  assign n3344 = n3343 & n3341;
  assign n3346 = {n3317, 1'b1};
  assign n3347 = n3346[0]; // extract
  assign n3348 = n3323[2]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3349 = n3344 ? n3347 : n3348;
  assign n3350 = n3346[1]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3351 = n3344 ? n3350 : n3317;
  assign n3352 = {n3351, n3349};
  assign n3353 = {n3337, n3335};
  assign n3354 = n3323[1:0]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3355 = n3325 ? n3353 : n3354;
  assign n3356 = n3352[0]; // extract
  assign n3357 = n3323[2]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3358 = n3325 ? n3357 : n3356;
  assign n3359 = n3352[1]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3360 = n3325 ? n3339 : n3359;
  /* TG68K_FPU.vhd:2473:63  */
  assign n3364 = ea_mode == 3'b000;
  /* TG68K_FPU.vhd:2475:74  */
  assign n3366 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:550:33  */
  assign n3373 = alu_operand_b[79]; // extract
  /* TG68K_FPU.vhd:551:37  */
  assign n3375 = alu_operand_b[78:64]; // extract
  /* TG68K_FPU.vhd:552:37  */
  assign n3377 = alu_operand_b[63:0]; // extract
  /* TG68K_FPU.vhd:558:29  */
  assign n3381 = n3375 == 15'b111111111111111;
  /* TG68K_FPU.vhd:560:36  */
  assign n3382 = alu_operand_b[63]; // extract
  /* TG68K_FPU.vhd:560:41  */
  assign n3383 = ~n3382;
  /* TG68K_FPU.vhd:560:58  */
  assign n3384 = alu_operand_b[62:0]; // extract
  /* TG68K_FPU.vhd:560:72  */
  assign n3386 = n3384 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:560:47  */
  assign n3387 = n3383 | n3386;
  assign n3390 = n3379[0]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3391 = n3387 ? 1'b1 : n3390;
  assign n3392 = n3379[1]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3393 = n3387 ? n3392 : 1'b1;
  assign n3394 = n3379[3]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3395 = n3387 ? n3394 : n3373;
  /* TG68K_FPU.vhd:568:32  */
  assign n3397 = n3375 == 15'b000000000000000;
  /* TG68K_FPU.vhd:568:68  */
  assign n3399 = n3377 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:568:55  */
  assign n3400 = n3399 & n3397;
  assign n3402 = {n3373, 1'b1};
  assign n3403 = n3402[0]; // extract
  assign n3404 = n3379[2]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3405 = n3400 ? n3403 : n3404;
  assign n3406 = n3402[1]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3407 = n3400 ? n3406 : n3373;
  assign n3408 = {n3407, n3405};
  assign n3409 = {n3393, n3391};
  assign n3410 = n3379[1:0]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3411 = n3381 ? n3409 : n3410;
  assign n3412 = n3408[0]; // extract
  assign n3413 = n3379[2]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3414 = n3381 ? n3413 : n3412;
  assign n3415 = n3408[1]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3416 = n3381 ? n3395 : n3415;
  /* TG68K_FPU.vhd:2481:77  */
  assign n3420 = fpu_operation == 7'b0001110;
  /* TG68K_FPU.vhd:2481:104  */
  assign n3422 = fpu_operation == 7'b0011101;
  /* TG68K_FPU.vhd:2481:87  */
  assign n3423 = n3420 | n3422;
  /* TG68K_FPU.vhd:2481:131  */
  assign n3425 = fpu_operation == 7'b0001111;
  /* TG68K_FPU.vhd:2481:114  */
  assign n3426 = n3423 | n3425;
  /* TG68K_FPU.vhd:2482:74  */
  assign n3428 = fpu_operation == 7'b0001100;
  /* TG68K_FPU.vhd:2481:141  */
  assign n3429 = n3426 | n3428;
  /* TG68K_FPU.vhd:2482:102  */
  assign n3431 = fpu_operation == 7'b0011100;
  /* TG68K_FPU.vhd:2482:85  */
  assign n3432 = n3429 | n3431;
  /* TG68K_FPU.vhd:2482:130  */
  assign n3434 = fpu_operation == 7'b0001010;
  /* TG68K_FPU.vhd:2482:113  */
  assign n3435 = n3432 | n3434;
  /* TG68K_FPU.vhd:2483:74  */
  assign n3437 = fpu_operation == 7'b0001011;
  /* TG68K_FPU.vhd:2482:141  */
  assign n3438 = n3435 | n3437;
  /* TG68K_FPU.vhd:2483:102  */
  assign n3440 = fpu_operation == 7'b0011001;
  /* TG68K_FPU.vhd:2483:85  */
  assign n3441 = n3438 | n3440;
  /* TG68K_FPU.vhd:2483:130  */
  assign n3443 = fpu_operation == 7'b0001001;
  /* TG68K_FPU.vhd:2483:113  */
  assign n3444 = n3441 | n3443;
  /* TG68K_FPU.vhd:2484:74  */
  assign n3446 = fpu_operation == 7'b0001101;
  /* TG68K_FPU.vhd:2483:141  */
  assign n3447 = n3444 | n3446;
  /* TG68K_FPU.vhd:2484:103  */
  assign n3449 = fpu_operation == 7'b0010000;
  /* TG68K_FPU.vhd:2484:86  */
  assign n3450 = n3447 | n3449;
  /* TG68K_FPU.vhd:2484:131  */
  assign n3452 = fpu_operation == 7'b0000111;
  /* TG68K_FPU.vhd:2484:114  */
  assign n3453 = n3450 | n3452;
  /* TG68K_FPU.vhd:2485:74  */
  assign n3455 = fpu_operation == 7'b0010001;
  /* TG68K_FPU.vhd:2484:144  */
  assign n3456 = n3453 | n3455;
  /* TG68K_FPU.vhd:2485:104  */
  assign n3458 = fpu_operation == 7'b0010010;
  /* TG68K_FPU.vhd:2485:87  */
  assign n3459 = n3456 | n3458;
  /* TG68K_FPU.vhd:2485:134  */
  assign n3461 = fpu_operation == 7'b0010100;
  /* TG68K_FPU.vhd:2485:117  */
  assign n3462 = n3459 | n3461;
  /* TG68K_FPU.vhd:2486:74  */
  assign n3464 = fpu_operation == 7'b0000101;
  /* TG68K_FPU.vhd:2485:145  */
  assign n3465 = n3462 | n3464;
  /* TG68K_FPU.vhd:2486:104  */
  assign n3467 = fpu_operation == 7'b0010101;
  /* TG68K_FPU.vhd:2486:87  */
  assign n3468 = n3465 | n3467;
  /* TG68K_FPU.vhd:2487:74  */
  assign n3470 = fpu_operation == 7'b0010110;
  /* TG68K_FPU.vhd:2486:116  */
  assign n3471 = n3468 | n3470;
  /* TG68K_FPU.vhd:2487:102  */
  assign n3473 = fpu_operation == 7'b0110000;
  /* TG68K_FPU.vhd:2487:85  */
  assign n3474 = n3471 | n3473;
  /* TG68K_FPU.vhd:2489:81  */
  assign n3475 = alu_operand_a[78:64]; // extract
  /* TG68K_FPU.vhd:2489:96  */
  assign n3477 = n3475 == 15'b111111111111111;
  /* TG68K_FPU.vhd:2491:89  */
  assign n3478 = alu_operand_a[63]; // extract
  /* TG68K_FPU.vhd:2491:117  */
  assign n3479 = alu_operand_a[62:0]; // extract
  /* TG68K_FPU.vhd:2491:131  */
  assign n3481 = n3479 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:2491:100  */
  assign n3482 = n3481 & n3478;
  /* TG68K_FPU.vhd:2495:92  */
  assign n3483 = alu_operand_a[63]; // extract
  /* TG68K_FPU.vhd:2495:120  */
  assign n3484 = alu_operand_a[62:0]; // extract
  /* TG68K_FPU.vhd:2495:134  */
  assign n3486 = n3484 == 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:2495:103  */
  assign n3487 = n3486 & n3483;
  /* TG68K_FPU.vhd:2498:89  */
  assign n3489 = fpu_operation == 7'b0001110;
  /* TG68K_FPU.vhd:2498:102  */
  assign n3491 = fpu_operation == 7'b0011101;
  /* TG68K_FPU.vhd:2498:102  */
  assign n3492 = n3489 | n3491;
  /* TG68K_FPU.vhd:2498:112  */
  assign n3494 = fpu_operation == 7'b0110000;
  /* TG68K_FPU.vhd:2498:112  */
  assign n3495 = n3492 | n3494;
  /* TG68K_FPU.vhd:2504:113  */
  assign n3496 = alu_operand_a[79]; // extract
  /* TG68K_FPU.vhd:2504:118  */
  assign n3497 = ~n3496;
  /* TG68K_FPU.vhd:2504:97  */
  assign n3499 = n3497 ? alu_operand_a : 80'b01111111111111111000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:2502:89  */
  assign n3501 = fpu_operation == 7'b0010100;
  /* TG68K_FPU.vhd:2502:103  */
  assign n3503 = fpu_operation == 7'b0010101;
  /* TG68K_FPU.vhd:2502:103  */
  assign n3504 = n3501 | n3503;
  /* TG68K_FPU.vhd:2502:115  */
  assign n3506 = fpu_operation == 7'b0010110;
  /* TG68K_FPU.vhd:2502:115  */
  assign n3507 = n3504 | n3506;
  assign n3508 = {n3507, n3495};
  /* TG68K_FPU.vhd:2497:81  */
  always @*
    case (n3508)
      2'b10: n3510 = n3298;
      2'b01: n3510 = n3298;
      default: n3510 = 4'b0101;
    endcase
  /* TG68K_FPU.vhd:2497:81  */
  always @*
    case (n3508)
      2'b10: n3512 = trans_start_operation;
      2'b01: n3512 = trans_start_operation;
      default: n3512 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:2497:81  */
  always @*
    case (n3508)
      2'b10: n3513 = trans_operation_code;
      2'b01: n3513 = trans_operation_code;
      default: n3513 = fpu_operation;
    endcase
  /* TG68K_FPU.vhd:2497:81  */
  always @*
    case (n3508)
      2'b10: n3514 = trans_operand;
      2'b01: n3514 = trans_operand;
      default: n3514 = alu_operand_a;
    endcase
  /* TG68K_FPU.vhd:2497:81  */
  always @*
    case (n3508)
      2'b10: n3516 = n3499;
      2'b01: n3516 = 80'b01111111111111111000000000000000000000000000000000000000000000000000000000000000;
      default: n3516 = result_data;
    endcase
  /* TG68K_FPU.vhd:2495:73  */
  assign n3518 = n3487 ? n3510 : 4'b0101;
  /* TG68K_FPU.vhd:2495:73  */
  assign n3520 = n3487 ? n3512 : 1'b1;
  /* TG68K_FPU.vhd:2495:73  */
  assign n3521 = n3487 ? n3513 : fpu_operation;
  /* TG68K_FPU.vhd:2495:73  */
  assign n3522 = n3487 ? n3514 : alu_operand_a;
  /* TG68K_FPU.vhd:2495:73  */
  assign n3523 = n3487 ? n3516 : result_data;
  /* TG68K_FPU.vhd:2491:73  */
  assign n3525 = n3482 ? 4'b0110 : n3518;
  /* TG68K_FPU.vhd:2491:73  */
  assign n3526 = n3482 ? trans_start_operation : n3520;
  /* TG68K_FPU.vhd:2491:73  */
  assign n3527 = n3482 ? trans_operation_code : n3521;
  /* TG68K_FPU.vhd:2491:73  */
  assign n3528 = n3482 ? trans_operand : n3522;
  /* TG68K_FPU.vhd:2491:73  */
  assign n3529 = n3482 ? alu_operand_a : n3523;
  /* TG68K_FPU.vhd:2529:107  */
  assign n3530 = fpcr_precision_valid & fpcr_rounding_mode_valid;
  /* TG68K_FPU.vhd:2535:88  */
  assign n3531 = fpcr[11]; // extract
  /* TG68K_FPU.vhd:2535:81  */
  assign n3533 = n3531 ? 1'b1 : n2926;
  /* TG68K_FPU.vhd:2535:81  */
  assign n3536 = n3531 ? 4'b1000 : 4'b0101;
  /* TG68K_FPU.vhd:2535:81  */
  assign n3538 = n3531 ? 8'b00010011 : n2930;
  /* TG68K_FPU.vhd:2535:81  */
  assign n3540 = n3531 ? trans_start_operation : 1'b1;
  /* TG68K_FPU.vhd:2529:73  */
  assign n3541 = n3530 ? n2926 : n3533;
  /* TG68K_FPU.vhd:2529:73  */
  assign n3543 = n3530 ? 4'b0101 : n3536;
  /* TG68K_FPU.vhd:2529:73  */
  assign n3544 = n3530 ? n2930 : n3538;
  /* TG68K_FPU.vhd:2529:73  */
  assign n3546 = n3530 ? 1'b1 : n3540;
  /* TG68K_FPU.vhd:2489:65  */
  assign n3547 = n3477 ? n2926 : n3541;
  /* TG68K_FPU.vhd:2489:65  */
  assign n3548 = n3477 ? n3525 : n3543;
  /* TG68K_FPU.vhd:2489:65  */
  assign n3549 = n3477 ? n2930 : n3544;
  /* TG68K_FPU.vhd:2489:65  */
  assign n3550 = n3477 ? n3526 : n3546;
  /* TG68K_FPU.vhd:2489:65  */
  assign n3551 = n3477 ? n3527 : fpu_operation;
  /* TG68K_FPU.vhd:2489:65  */
  assign n3552 = n3477 ? n3528 : alu_operand_a;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3553 = n3575 ? n3529 : result_data;
  /* TG68K_FPU.vhd:2552:99  */
  assign n3554 = fpcr_precision_valid & fpcr_rounding_mode_valid;
  /* TG68K_FPU.vhd:2560:80  */
  assign n3555 = fpcr[11]; // extract
  /* TG68K_FPU.vhd:2560:73  */
  assign n3557 = n3555 ? 1'b1 : n2926;
  /* TG68K_FPU.vhd:2560:73  */
  assign n3561 = n3555 ? 8'b00010011 : n2930;
  /* TG68K_FPU.vhd:2552:65  */
  assign n3562 = n3554 ? n2926 : n3557;
  /* TG68K_FPU.vhd:2552:65  */
  assign n3564 = n3554 ? n2930 : n3561;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3565 = n3474 ? n3547 : n3562;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3567 = n3474 ? n3548 : 4'b0101;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3568 = n3474 ? n3549 : n3564;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3570 = n3474 ? n3300 : 1'b1;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3571 = n3474 ? n3301 : fpu_operation;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3572 = n3474 ? n3550 : trans_start_operation;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3573 = n3474 ? n3551 : trans_operation_code;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3574 = n3474 ? n3552 : trans_operand;
  /* TG68K_FPU.vhd:2481:57  */
  assign n3575 = n3477 & n3474;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3576 = n3366 ? n2926 : n3565;
  assign n3577 = {n3416, n3414, n3411};
  assign n3578 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:2473:49  */
  assign n3579 = n3591 ? n3577 : n3578;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3581 = n3366 ? 4'b0111 : n3567;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3582 = n3366 ? n2930 : n3568;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3583 = n3366 ? n3300 : n3570;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3584 = n3366 ? n3301 : n3571;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3585 = n3366 ? trans_start_operation : n3572;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3586 = n3366 ? trans_operation_code : n3573;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3587 = n3366 ? trans_operand : n3574;
  /* TG68K_FPU.vhd:2475:57  */
  assign n3588 = n3366 ? result_data : n3553;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3589 = n3364 ? n3576 : n2926;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3591 = n3366 & n3364;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3592 = n3364 ? n3581 : n3298;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3593 = n3364 ? n3582 : n2930;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3594 = n3364 ? n3583 : n3300;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3595 = n3364 ? n3584 : n3301;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3596 = n3364 ? n3585 : trans_start_operation;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3597 = n3364 ? n3586 : trans_operation_code;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3598 = n3364 ? n3587 : trans_operand;
  /* TG68K_FPU.vhd:2473:49  */
  assign n3599 = n3364 ? n3588 : result_data;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3600 = n3310 ? n2926 : n3589;
  assign n3601 = {n3360, n3358, n3355};
  /* TG68K_FPU.vhd:2466:49  */
  assign n3602 = n3310 ? n3601 : n3579;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3604 = n3310 ? 4'b0111 : n3592;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3605 = n3310 ? n2930 : n3593;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3606 = n3310 ? n3300 : n3594;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3607 = n3310 ? n3301 : n3595;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3608 = n3310 ? trans_start_operation : n3596;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3609 = n3310 ? trans_operation_code : n3597;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3610 = n3310 ? trans_operand : n3598;
  /* TG68K_FPU.vhd:2466:49  */
  assign n3611 = n3310 ? result_data : n3599;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3612 = n2915 ? fpu_exception_i : n3600;
  assign n3613 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:2167:49  */
  assign n3614 = n2915 ? n3613 : n3602;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3615 = n2915 ? fpu_state : n3604;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3616 = n2915 ? exception_code_internal : n3605;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3618 = n2915 ? 1'b0 : n3606;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3619 = n2915 ? alu_operation_code : n3607;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3620 = n2915 ? alu_operand_a : n2931;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3621 = n2915 ? alu_operand_b : n3302;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3622 = n2915 ? trans_start_operation : n3608;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3623 = n2915 ? trans_operation_code : n3609;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3624 = n2915 ? trans_operand : n3610;
  /* TG68K_FPU.vhd:2167:49  */
  assign n3625 = n2915 ? result_data : n3611;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3626 = n2799 ? fpu_exception_i : n3612;
  assign n3627 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:2095:49  */
  assign n3628 = n2799 ? n3627 : n3614;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3630 = n2799 ? 4'b0101 : n3615;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3631 = n2799 ? exception_code_internal : n3616;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3633 = n2799 ? 1'b1 : n3618;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3635 = n2799 ? fpu_operation : n3619;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3636 = n2799 ? alu_operand_a : n3620;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3637 = n2799 ? n2910 : n3621;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3638 = n2799 ? trans_start_operation : n3622;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3639 = n2799 ? trans_operation_code : n3623;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3640 = n2799 ? trans_operand : n3624;
  /* TG68K_FPU.vhd:2095:49  */
  assign n3641 = n2799 ? result_data : n3625;
  /* TG68K_FPU.vhd:2088:41  */
  assign n3643 = fpu_state == 4'b0010;
  /* TG68K_FPU.vhd:2578:68  */
  assign n3644 = {24'b0, timeout_counter};  //  uext
  /* TG68K_FPU.vhd:2578:68  */
  assign n3646 = $signed(n3644) < $signed(32'b00000000000000000000000001000000);
  /* TG68K_FPU.vhd:2579:92  */
  assign n3647 = {24'b0, timeout_counter};  //  uext
  /* TG68K_FPU.vhd:2579:92  */
  assign n3649 = n3647 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:2579:76  */
  assign n3650 = n3649[7:0];  // trunc
  /* TG68K_FPU.vhd:2578:49  */
  assign n3651 = n3646 ? n3650 : timeout_counter;
  /* TG68K_FPU.vhd:2584:77  */
  assign n3652 = ~fpcr_rounding_mode_valid;
  /* TG68K_FPU.vhd:2591:64  */
  assign n3654 = fpcr[11]; // extract
  /* TG68K_FPU.vhd:2584:49  */
  assign n3656 = n3661 ? 1'b1 : fpu_exception_i;
  /* TG68K_FPU.vhd:2584:49  */
  assign n3658 = n3668 ? 4'b1000 : fpu_state;
  /* TG68K_FPU.vhd:2584:49  */
  assign n3660 = n3669 ? 8'b00010011 : exception_code_internal;
  /* TG68K_FPU.vhd:2584:49  */
  assign n3661 = n3654 & n3652;
  assign n3662 = fpcr[15:14]; // extract
  /* TG68K_FPU.vhd:2584:49  */
  assign n3663 = n3652 ? 2'b00 : n3662;
  /* TG68K_FPU.vhd:2584:49  */
  assign n3667 = n3652 ? 1'b1 : fpcr_rounding_mode_valid;
  /* TG68K_FPU.vhd:2584:49  */
  assign n3668 = n3654 & n3652;
  /* TG68K_FPU.vhd:2584:49  */
  assign n3669 = n3654 & n3652;
  /* TG68K_FPU.vhd:2599:73  */
  assign n3670 = ~fpcr_precision_valid;
  /* TG68K_FPU.vhd:2606:64  */
  assign n3672 = fpcr[11]; // extract
  /* TG68K_FPU.vhd:2599:49  */
  assign n3674 = n3679 ? 1'b1 : n3656;
  /* TG68K_FPU.vhd:2599:49  */
  assign n3676 = n3686 ? 4'b1000 : n3658;
  /* TG68K_FPU.vhd:2599:49  */
  assign n3678 = n3687 ? 8'b00010011 : n3660;
  /* TG68K_FPU.vhd:2599:49  */
  assign n3679 = n3672 & n3670;
  assign n3680 = fpcr[7:6]; // extract
  /* TG68K_FPU.vhd:2599:49  */
  assign n3681 = n3670 ? 2'b00 : n3680;
  /* TG68K_FPU.vhd:2599:49  */
  assign n3685 = n3670 ? 1'b1 : fpcr_precision_valid;
  /* TG68K_FPU.vhd:2599:49  */
  assign n3686 = n3672 & n3670;
  /* TG68K_FPU.vhd:2599:49  */
  assign n3687 = n3672 & n3670;
  /* TG68K_FPU.vhd:2614:66  */
  assign n3689 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:2614:96  */
  assign n3691 = decoder_ea_mode == 3'b000;
  /* TG68K_FPU.vhd:2614:76  */
  assign n3692 = n3691 & n3689;
  /* TG68K_FPU.vhd:2620:69  */
  assign n3694 = fpu_operation == 7'b1000000;
  /* TG68K_FPU.vhd:2626:76  */
  assign n3695 = {24'b0, timeout_counter};  //  uext
  /* TG68K_FPU.vhd:2626:76  */
  assign n3697 = $signed(n3695) > $signed(32'b00000000000000000000000010000000);
  /* TG68K_FPU.vhd:2620:49  */
  assign n3699 = n4010 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:2626:57  */
  assign n3701 = n3697 ? 4'b0000 : n3676;
  /* TG68K_FPU.vhd:2631:81  */
  assign n3702 = alu_operation_done | alu_result_valid;
  /* TG68K_FPU.vhd:2631:139  */
  assign n3703 = trans_operation_done | trans_result_valid;
  /* TG68K_FPU.vhd:2631:108  */
  assign n3704 = n3702 | n3703;
  /* TG68K_FPU.vhd:2636:87  */
  assign n3705 = trans_operation_done | trans_result_valid;
  /* TG68K_FPU.vhd:2636:57  */
  assign n3706 = n3705 ? trans_result : alu_result;
  /* TG68K_FPU.vhd:2636:57  */
  assign n3707 = n3705 ? trans_overflow : alu_overflow;
  /* TG68K_FPU.vhd:2636:57  */
  assign n3708 = n3705 ? trans_underflow : alu_underflow;
  /* TG68K_FPU.vhd:2636:57  */
  assign n3709 = n3705 ? trans_inexact : alu_inexact;
  /* TG68K_FPU.vhd:2636:57  */
  assign n3710 = n3705 ? trans_invalid : alu_invalid;
  /* TG68K_FPU.vhd:2656:75  */
  assign n3712 = fpu_operation == 7'b0100001;
  /* TG68K_FPU.vhd:2656:102  */
  assign n3714 = fpu_operation == 7'b0100101;
  /* TG68K_FPU.vhd:2656:85  */
  assign n3715 = n3712 | n3714;
  assign n3716 = exception_fpsr_out[23:16]; // extract
  /* TG68K_FPU.vhd:2656:57  */
  assign n3717 = n3715 ? alu_quotient_byte : n3716;
  assign n3718 = exception_fpsr_out[31:24]; // extract
  assign n3719 = exception_fpsr_out[15:0]; // extract
  /* TG68K_FPU.vhd:613:28  */
  assign n3730 = fpcr[7:6]; // extract
  /* TG68K_FPU.vhd:613:41  */
  assign n3732 = n3730 == 2'b11;
  /* TG68K_FPU.vhd:613:17  */
  assign n3736 = n3732 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:613:17  */
  assign n3742 = n3732 ? 1'b0 : 1'bX;
  /* TG68K_FPU.vhd:618:28  */
  assign n3743 = fpcr[31:16]; // extract
  /* TG68K_FPU.vhd:618:43  */
  assign n3745 = n3743 != 16'b0000000000000000;
  /* TG68K_FPU.vhd:618:65  */
  assign n3746 = fpcr[5:0]; // extract
  /* TG68K_FPU.vhd:618:78  */
  assign n3748 = n3746 != 6'b000000;
  /* TG68K_FPU.vhd:618:54  */
  assign n3749 = n3745 | n3748;
  /* TG68K_FPU.vhd:618:17  */
  assign n3752 = n3759 ? 1'b0 : n3736;
  /* TG68K_FPU.vhd:618:17  */
  assign n3755 = n3761 ? 1'b0 : n3742;
  /* TG68K_FPU.vhd:618:17  */
  assign n3756 = n3736 & n3749;
  /* TG68K_FPU.vhd:618:17  */
  assign n3758 = n3736 & n3749;
  /* TG68K_FPU.vhd:618:17  */
  assign n3759 = n3756 & n3736;
  /* TG68K_FPU.vhd:618:17  */
  assign n3761 = n3758 & n3736;
  /* TG68K_FPU.vhd:623:17  */
  assign n3767 = n3752 ? 1'b1 : n3755;
  /* TG68K_FPU.vhd:641:56  */
  assign n3768 = fpcr[7:6]; // extract
  /* TG68K_FPU.vhd:641:69  */
  assign n3770 = n3768 != 2'b11;
  /* TG68K_FPU.vhd:641:44  */
  assign n3771 = n3770 & n3767;
  /* TG68K_FPU.vhd:642:40  */
  assign n3772 = fpcr[7:6]; // extract
  /* TG68K_FPU.vhd:641:17  */
  assign n3774 = n3771 ? n3772 : 2'b00;
  /* TG68K_FPU.vhd:2675:81  */
  assign n3776 = fpcr_precision_bits == 2'b00;
  /* TG68K_FPU.vhd:2681:104  */
  assign n3777 = final_result[78:64]; // extract
  /* TG68K_FPU.vhd:2681:119  */
  assign n3779 = n3777 == 15'b000000000000000;
  /* TG68K_FPU.vhd:2684:107  */
  assign n3780 = final_result[78:64]; // extract
  /* TG68K_FPU.vhd:2684:122  */
  assign n3782 = n3780 == 15'b111111111111111;
  /* TG68K_FPU.vhd:2690:124  */
  assign n3783 = final_result[79]; // extract
  /* TG68K_FPU.vhd:2690:129  */
  assign n3785 = {n3783, 15'b011111111111111};
  /* TG68K_FPU.vhd:2690:149  */
  assign n3787 = {n3785, 1'b1};
  /* TG68K_FPU.vhd:2690:169  */
  assign n3788 = final_result[62:40]; // extract
  /* TG68K_FPU.vhd:2690:155  */
  assign n3789 = {n3787, n3788};
  /* TG68K_FPU.vhd:2690:184  */
  assign n3791 = {n3789, 40'b0000000000000000000000000000000000000000};
  /* TG68K_FPU.vhd:2684:89  */
  assign n3792 = n3782 ? final_result : n3791;
  /* TG68K_FPU.vhd:2681:89  */
  assign n3794 = n3779 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3792;
  /* TG68K_FPU.vhd:2677:81  */
  assign n3796 = fpcr_precision_bits == 2'b01;
  /* TG68K_FPU.vhd:2695:104  */
  assign n3797 = final_result[78:64]; // extract
  /* TG68K_FPU.vhd:2695:119  */
  assign n3799 = n3797 == 15'b000000000000000;
  /* TG68K_FPU.vhd:2698:107  */
  assign n3800 = final_result[78:64]; // extract
  /* TG68K_FPU.vhd:2698:122  */
  assign n3802 = n3800 == 15'b111111111111111;
  /* TG68K_FPU.vhd:2704:124  */
  assign n3803 = final_result[79]; // extract
  /* TG68K_FPU.vhd:2704:129  */
  assign n3805 = {n3803, 15'b011111111111111};
  /* TG68K_FPU.vhd:2704:163  */
  assign n3806 = final_result[63:0]; // extract
  /* TG68K_FPU.vhd:2704:149  */
  assign n3807 = {n3805, n3806};
  /* TG68K_FPU.vhd:2698:89  */
  assign n3808 = n3802 ? final_result : n3807;
  /* TG68K_FPU.vhd:2695:89  */
  assign n3810 = n3799 ? 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000 : n3808;
  /* TG68K_FPU.vhd:2692:81  */
  assign n3812 = fpcr_precision_bits == 2'b10;
  assign n3813 = {n3812, n3796, n3776};
  /* TG68K_FPU.vhd:2674:73  */
  always @*
    case (n3813)
      3'b100: n3815 = n3685;
      3'b010: n3815 = n3685;
      3'b001: n3815 = n3685;
      default: n3815 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:2674:73  */
  always @*
    case (n3813)
      3'b100: n3816 = n3810;
      3'b010: n3816 = n3794;
      3'b001: n3816 = final_result;
      default: n3816 = final_result;
    endcase
  /* TG68K_FPU.vhd:2671:65  */
  assign n3817 = fpcr_precision_valid ? n3815 : n3685;
  /* TG68K_FPU.vhd:2671:65  */
  assign n3818 = fpcr_precision_valid ? n3774 : fpcr_precision_bits;
  /* TG68K_FPU.vhd:2671:65  */
  assign n3819 = fpcr_precision_valid ? n3816 : final_result;
  /* TG68K_FPU.vhd:2661:57  */
  assign n3821 = exception_pending_internal ? 1'b1 : n3674;
  /* TG68K_FPU.vhd:2661:57  */
  assign n3822 = exception_pending_internal ? n3685 : n3817;
  /* TG68K_FPU.vhd:2661:57  */
  assign n3823 = exception_pending_internal ? fpcr_precision_bits : n3818;
  /* TG68K_FPU.vhd:2661:57  */
  assign n3826 = exception_pending_internal ? 4'b1000 : 4'b0110;
  /* TG68K_FPU.vhd:2661:57  */
  assign n3827 = exception_pending_internal ? exception_vector_internal : n3678;
  /* TG68K_FPU.vhd:2661:57  */
  assign n3828 = exception_pending_internal ? exception_corrected_result : n3819;
  /* TG68K_FPU.vhd:2719:71  */
  assign n3829 = {24'b0, timeout_counter};  //  uext
  /* TG68K_FPU.vhd:2719:71  */
  assign n3831 = $signed(n3829) >= $signed(32'b00000000000000000000000001000000);
  /* TG68K_FPU.vhd:2722:74  */
  assign n3833 = fpu_operation == 7'b0000000;
  /* TG68K_FPU.vhd:2722:102  */
  assign n3835 = fpu_operation == 7'b0011000;
  /* TG68K_FPU.vhd:2722:85  */
  assign n3836 = n3833 | n3835;
  /* TG68K_FPU.vhd:2722:129  */
  assign n3838 = fpu_operation == 7'b0011010;
  /* TG68K_FPU.vhd:2722:112  */
  assign n3839 = n3836 | n3838;
  /* TG68K_FPU.vhd:2724:82  */
  assign n3841 = fpu_operation == 7'b0000000;
  /* TG68K_FPU.vhd:2726:85  */
  assign n3843 = fpu_operation == 7'b0011000;
  /* TG68K_FPU.vhd:2727:107  */
  assign n3844 = alu_operand_a[78:0]; // extract
  /* TG68K_FPU.vhd:2727:92  */
  assign n3846 = {1'b0, n3844};
  /* TG68K_FPU.vhd:2728:85  */
  assign n3848 = fpu_operation == 7'b0011010;
  /* TG68K_FPU.vhd:2729:106  */
  assign n3849 = alu_operand_a[79]; // extract
  /* TG68K_FPU.vhd:2729:89  */
  assign n3850 = ~n3849;
  /* TG68K_FPU.vhd:2729:127  */
  assign n3851 = alu_operand_a[78:0]; // extract
  /* TG68K_FPU.vhd:2729:112  */
  assign n3852 = {n3850, n3851};
  /* TG68K_FPU.vhd:2728:65  */
  assign n3853 = n3848 ? n3852 : result_data;
  /* TG68K_FPU.vhd:2726:65  */
  assign n3854 = n3843 ? n3846 : n3853;
  /* TG68K_FPU.vhd:2724:65  */
  assign n3855 = n3841 ? alu_operand_b : n3854;
  /* TG68K_FPU.vhd:2732:77  */
  assign n3857 = fpu_operation == 7'b0111010;
  /* TG68K_FPU.vhd:2735:76  */
  assign n3859 = ea_mode == 3'b000;
  /* TG68K_FPU.vhd:550:33  */
  assign n3866 = alu_operand_b[79]; // extract
  /* TG68K_FPU.vhd:551:37  */
  assign n3868 = alu_operand_b[78:64]; // extract
  /* TG68K_FPU.vhd:552:37  */
  assign n3870 = alu_operand_b[63:0]; // extract
  /* TG68K_FPU.vhd:558:29  */
  assign n3874 = n3868 == 15'b111111111111111;
  /* TG68K_FPU.vhd:560:36  */
  assign n3875 = alu_operand_b[63]; // extract
  /* TG68K_FPU.vhd:560:41  */
  assign n3876 = ~n3875;
  /* TG68K_FPU.vhd:560:58  */
  assign n3877 = alu_operand_b[62:0]; // extract
  /* TG68K_FPU.vhd:560:72  */
  assign n3879 = n3877 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:560:47  */
  assign n3880 = n3876 | n3879;
  assign n3883 = n3872[0]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3884 = n3880 ? 1'b1 : n3883;
  assign n3885 = n3872[1]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3886 = n3880 ? n3885 : 1'b1;
  assign n3887 = n3872[3]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3888 = n3880 ? n3887 : n3866;
  /* TG68K_FPU.vhd:568:32  */
  assign n3890 = n3868 == 15'b000000000000000;
  /* TG68K_FPU.vhd:568:68  */
  assign n3892 = n3870 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:568:55  */
  assign n3893 = n3892 & n3890;
  assign n3895 = {n3866, 1'b1};
  assign n3896 = n3895[0]; // extract
  assign n3897 = n3872[2]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3898 = n3893 ? n3896 : n3897;
  assign n3899 = n3895[1]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3900 = n3893 ? n3899 : n3866;
  assign n3901 = {n3900, n3898};
  assign n3902 = {n3886, n3884};
  assign n3903 = n3872[1:0]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3904 = n3874 ? n3902 : n3903;
  assign n3905 = n3901[0]; // extract
  assign n3906 = n3872[2]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3907 = n3874 ? n3906 : n3905;
  assign n3908 = n3901[1]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3909 = n3874 ? n3888 : n3908;
  /* TG68K_FPU.vhd:550:33  */
  assign n3918 = alu_operand_a[79]; // extract
  /* TG68K_FPU.vhd:551:37  */
  assign n3920 = alu_operand_a[78:64]; // extract
  /* TG68K_FPU.vhd:552:37  */
  assign n3922 = alu_operand_a[63:0]; // extract
  /* TG68K_FPU.vhd:558:29  */
  assign n3926 = n3920 == 15'b111111111111111;
  /* TG68K_FPU.vhd:560:36  */
  assign n3927 = alu_operand_a[63]; // extract
  /* TG68K_FPU.vhd:560:41  */
  assign n3928 = ~n3927;
  /* TG68K_FPU.vhd:560:58  */
  assign n3929 = alu_operand_a[62:0]; // extract
  /* TG68K_FPU.vhd:560:72  */
  assign n3931 = n3929 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:560:47  */
  assign n3932 = n3928 | n3931;
  assign n3935 = n3924[0]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3936 = n3932 ? 1'b1 : n3935;
  assign n3937 = n3924[1]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3938 = n3932 ? n3937 : 1'b1;
  assign n3939 = n3924[3]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n3940 = n3932 ? n3939 : n3918;
  /* TG68K_FPU.vhd:568:32  */
  assign n3942 = n3920 == 15'b000000000000000;
  /* TG68K_FPU.vhd:568:68  */
  assign n3944 = n3922 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:568:55  */
  assign n3945 = n3944 & n3942;
  assign n3947 = {n3918, 1'b1};
  assign n3948 = n3947[0]; // extract
  assign n3949 = n3924[2]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3950 = n3945 ? n3948 : n3949;
  assign n3951 = n3947[1]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n3952 = n3945 ? n3951 : n3918;
  assign n3953 = {n3952, n3950};
  assign n3954 = {n3938, n3936};
  assign n3955 = n3924[1:0]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3956 = n3926 ? n3954 : n3955;
  assign n3957 = n3953[0]; // extract
  assign n3958 = n3924[2]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3959 = n3926 ? n3958 : n3957;
  assign n3960 = n3953[1]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n3961 = n3926 ? n3940 : n3960;
  assign n3964 = {n3961, n3959, n3956};
  assign n3965 = {n3909, n3907, n3904};
  /* TG68K_FPU.vhd:2735:65  */
  assign n3966 = n3859 ? n3965 : n3964;
  /* TG68K_FPU.vhd:2732:57  */
  assign n3968 = n3857 ? n3674 : 1'b1;
  assign n3969 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:2732:57  */
  assign n3970 = n3857 ? n3966 : n3969;
  /* TG68K_FPU.vhd:2732:57  */
  assign n3973 = n3857 ? 4'b0111 : 4'b1000;
  /* TG68K_FPU.vhd:2732:57  */
  assign n3975 = n3857 ? n3678 : 8'b00001011;
  /* TG68K_FPU.vhd:2722:57  */
  assign n3976 = n3839 ? n3674 : n3968;
  assign n3977 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:2722:57  */
  assign n3978 = n3839 ? n3977 : n3970;
  /* TG68K_FPU.vhd:2722:57  */
  assign n3980 = n3839 ? 4'b0110 : n3973;
  /* TG68K_FPU.vhd:2722:57  */
  assign n3981 = n3839 ? n3678 : n3975;
  /* TG68K_FPU.vhd:2719:49  */
  assign n3982 = n3990 ? n3855 : result_data;
  /* TG68K_FPU.vhd:2719:49  */
  assign n3983 = n3831 ? n3976 : n3674;
  assign n3984 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:2719:49  */
  assign n3985 = n3831 ? n3978 : n3984;
  /* TG68K_FPU.vhd:2719:49  */
  assign n3986 = n3831 ? n3980 : n3676;
  /* TG68K_FPU.vhd:2719:49  */
  assign n3988 = n3831 ? 8'b00000000 : n3651;
  /* TG68K_FPU.vhd:2719:49  */
  assign n3989 = n3831 ? n3981 : n3678;
  /* TG68K_FPU.vhd:2719:49  */
  assign n3990 = n3839 & n3831;
  /* TG68K_FPU.vhd:2631:49  */
  assign n3991 = n3704 ? n3821 : n3983;
  assign n3992 = {n3718, n3717, n3719};
  assign n3993 = n3992[27:0]; // extract
  assign n3994 = fpsr[27:0]; // extract
  /* TG68K_FPU.vhd:2631:49  */
  assign n3995 = n3704 ? n3993 : n3994;
  assign n3996 = n3992[31:28]; // extract
  /* TG68K_FPU.vhd:2631:49  */
  assign n3997 = n3704 ? n3996 : n3985;
  /* TG68K_FPU.vhd:2631:49  */
  assign n3998 = n3704 ? n3822 : n3685;
  /* TG68K_FPU.vhd:2631:49  */
  assign n3999 = n3704 ? n3823 : fpcr_precision_bits;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4000 = n3704 ? n3826 : n3986;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4002 = n3704 ? 8'b00000000 : n3988;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4003 = n3704 ? n3827 : n3989;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4004 = n3704 ? n3706 : final_result;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4005 = n3704 ? n3707 : final_overflow;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4006 = n3704 ? n3708 : final_underflow;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4007 = n3704 ? n3709 : final_inexact;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4008 = n3704 ? n3710 : final_invalid;
  /* TG68K_FPU.vhd:2631:49  */
  assign n4009 = n3704 ? n3828 : n3982;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4010 = n3697 & n3694;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4011 = n3694 ? n3674 : n3991;
  assign n4012 = {n3997, n3995};
  /* TG68K_FPU.vhd:2620:49  */
  assign n4013 = n3694 ? fpsr : n4012;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4014 = n3694 ? n3685 : n3998;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4015 = n3694 ? fpcr_precision_bits : n3999;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4016 = n3694 ? n3701 : n4000;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4017 = n3694 ? n3651 : n4002;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4018 = n3694 ? n3678 : n4003;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4019 = n3694 ? final_result : n4004;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4020 = n3694 ? final_overflow : n4005;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4021 = n3694 ? final_underflow : n4006;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4022 = n3694 ? final_inexact : n4007;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4023 = n3694 ? final_invalid : n4008;
  /* TG68K_FPU.vhd:2620:49  */
  assign n4024 = n3694 ? result_data : n4009;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4026 = n3692 ? 1'b1 : n3699;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4027 = n3692 ? n3674 : n4011;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4028 = n3692 ? fpsr : n4013;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4029 = n3692 ? n3685 : n4014;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4030 = n3692 ? fpcr_precision_bits : n4015;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4032 = n3692 ? 4'b0000 : n4016;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4034 = n3692 ? 8'b00000000 : n4017;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4035 = n3692 ? n3678 : n4018;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4036 = n3692 ? final_result : n4019;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4037 = n3692 ? final_overflow : n4020;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4038 = n3692 ? final_underflow : n4021;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4039 = n3692 ? final_inexact : n4022;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4040 = n3692 ? final_invalid : n4023;
  /* TG68K_FPU.vhd:2614:49  */
  assign n4041 = n3692 ? result_data : n4024;
  /* TG68K_FPU.vhd:2573:41  */
  assign n4043 = fpu_state == 4'b0101;
  /* TG68K_FPU.vhd:2755:41  */
  assign n4045 = fpu_state == 4'b0011;
  /* TG68K_FPU.vhd:2759:41  */
  assign n4047 = fpu_state == 4'b0100;
  /* TG68K_FPU.vhd:2766:66  */
  assign n4049 = fpu_operation == 7'b1000001;
  /* TG68K_FPU.vhd:2770:68  */
  assign n4050 = {28'b0, dest_reg};  //  uext
  /* TG68K_FPU.vhd:2770:99  */
  assign n4051 = {1'b0, n4050};  //  uext
  /* TG68K_FPU.vhd:2770:99  */
  assign n4053 = $signed(n4051) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:2770:65  */
  assign n4055 = n4053 ? fpu_exception_i : 1'b1;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4057 = n4069 ? 1'b1 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4058 = n4070 ? dest_reg : fp_reg_write_addr;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4059 = n4071 ? constrom_result : fp_reg_write_data;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4061 = n4072 ? 1'b1 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:2770:65  */
  assign n4065 = n4053 ? exception_code_internal : 8'b00010100;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4067 = constrom_valid ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4068 = n4330 ? n4055 : fpu_exception_i;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4069 = n4053 & constrom_valid;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4070 = n4053 & constrom_valid;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4071 = n4053 & constrom_valid;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4072 = n4053 & constrom_valid;
  /* TG68K_FPU.vhd:2768:57  */
  assign n4074 = constrom_valid ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4075 = n4345 ? n4065 : exception_code_internal;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4077 = n4346 ? 1'b0 : rom_read_enable;
  /* TG68K_FPU.vhd:2788:74  */
  assign n4079 = fpu_operation == 7'b0110000;
  /* TG68K_FPU.vhd:2791:68  */
  assign n4080 = {28'b0, dest_reg};  //  uext
  /* TG68K_FPU.vhd:2791:99  */
  assign n4081 = {1'b0, n4080};  //  uext
  /* TG68K_FPU.vhd:2791:99  */
  assign n4083 = $signed(n4081) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:2791:65  */
  assign n4091 = n4083 ? 1'b1 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:2791:65  */
  assign n4092 = n4083 ? dest_reg : fp_reg_write_addr;
  /* TG68K_FPU.vhd:2791:65  */
  assign n4093 = n4083 ? result_data : fp_reg_write_data;
  /* TG68K_FPU.vhd:2791:65  */
  assign n4095 = n4083 ? 1'b1 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:2803:102  */
  assign n4096 = extension_word[2:0]; // extract
  /* TG68K_FPU.vhd:2803:68  */
  assign n4097 = {28'b0, n4096};  //  uext
  /* TG68K_FPU.vhd:2803:117  */
  assign n4098 = {1'b0, n4097};  //  uext
  /* TG68K_FPU.vhd:2803:117  */
  assign n4100 = $signed(n4098) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:2804:87  */
  assign n4101 = result_data[78:64]; // extract
  /* TG68K_FPU.vhd:2804:102  */
  assign n4103 = n4101 == 15'b111111111111111;
  /* TG68K_FPU.vhd:2807:116  */
  assign n4104 = extension_word[2:0]; // extract
  /* TG68K_FPU.vhd:2818:97  */
  assign n4111 = alu_operand_a[78:64]; // extract
  /* TG68K_FPU.vhd:2818:112  */
  assign n4113 = $unsigned(n4111) < $unsigned(15'b100000000000001);
  /* TG68K_FPU.vhd:2821:124  */
  assign n4114 = extension_word[2:0]; // extract
  /* TG68K_FPU.vhd:2828:100  */
  assign n4121 = alu_operand_a[78:64]; // extract
  /* TG68K_FPU.vhd:2828:115  */
  assign n4123 = $unsigned(n4121) > $unsigned(15'b100000000010100);
  /* TG68K_FPU.vhd:2831:124  */
  assign n4124 = extension_word[2:0]; // extract
  /* TG68K_FPU.vhd:2842:105  */
  assign n4131 = alu_operand_a[78:64]; // extract
  /* TG68K_FPU.vhd:2842:120  */
  assign n4133 = n4131 == 15'b100000000000000;
  /* TG68K_FPU.vhd:2845:132  */
  assign n4134 = extension_word[2:0]; // extract
  /* TG68K_FPU.vhd:2852:108  */
  assign n4141 = alu_operand_a[78:64]; // extract
  /* TG68K_FPU.vhd:2852:123  */
  assign n4143 = n4141 == 15'b100000000000001;
  /* TG68K_FPU.vhd:2855:132  */
  assign n4144 = extension_word[2:0]; // extract
  /* TG68K_FPU.vhd:2866:132  */
  assign n4151 = extension_word[2:0]; // extract
  /* TG68K_FPU.vhd:2852:89  */
  assign n4160 = n4143 ? n4144 : n4151;
  /* TG68K_FPU.vhd:2852:89  */
  assign n4163 = n4143 ? 80'b10111111111111101101010100101100110101000100110011101000101000000000000000000000 : 80'b00111111111111110000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:2842:89  */
  assign n4166 = n4133 ? n4134 : n4160;
  /* TG68K_FPU.vhd:2842:89  */
  assign n4168 = n4133 ? 80'b00111111111111101000101001010001010000000111110110100111001111111000000000000000 : n4163;
  /* TG68K_FPU.vhd:2828:81  */
  assign n4171 = n4123 ? n4124 : n4166;
  /* TG68K_FPU.vhd:2828:81  */
  assign n4173 = n4123 ? 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000 : n4168;
  /* TG68K_FPU.vhd:2818:81  */
  assign n4176 = n4113 ? n4114 : n4171;
  /* TG68K_FPU.vhd:2818:81  */
  assign n4178 = n4113 ? 80'b00111111111111111000000000000000000000000000000000000000000000000000000000000000 : n4173;
  /* TG68K_FPU.vhd:2804:73  */
  assign n4181 = n4103 ? n4104 : n4176;
  /* TG68K_FPU.vhd:2804:73  */
  assign n4182 = n4103 ? result_data : n4178;
  /* TG68K_FPU.vhd:2803:65  */
  assign n4186 = n4100 ? 1'b1 : n4091;
  /* TG68K_FPU.vhd:2803:65  */
  assign n4187 = n4100 ? n4181 : n4092;
  /* TG68K_FPU.vhd:2803:65  */
  assign n4188 = n4100 ? n4182 : n4093;
  /* TG68K_FPU.vhd:2803:65  */
  assign n4190 = n4100 ? 1'b1 : n4095;
  /* TG68K_FPU.vhd:2877:77  */
  assign n4192 = fpu_operation != 7'b0111010;
  /* TG68K_FPU.vhd:2877:106  */
  assign n4194 = fpu_operation != 7'b0111000;
  /* TG68K_FPU.vhd:2877:88  */
  assign n4195 = n4194 & n4192;
  /* TG68K_FPU.vhd:2880:68  */
  assign n4196 = {28'b0, dest_reg};  //  uext
  /* TG68K_FPU.vhd:2880:99  */
  assign n4197 = {1'b0, n4196};  //  uext
  /* TG68K_FPU.vhd:2880:99  */
  assign n4199 = $signed(n4197) <= $signed(32'b00000000000000000000000000000111);
  /* TG68K_FPU.vhd:2877:57  */
  assign n4207 = n4214 ? 1'b1 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:2877:57  */
  assign n4208 = n4215 ? dest_reg : fp_reg_write_addr;
  /* TG68K_FPU.vhd:2877:57  */
  assign n4209 = n4216 ? result_data : fp_reg_write_data;
  /* TG68K_FPU.vhd:2877:57  */
  assign n4211 = n4217 ? 1'b1 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:2877:57  */
  assign n4214 = n4199 & n4195;
  /* TG68K_FPU.vhd:2877:57  */
  assign n4215 = n4199 & n4195;
  /* TG68K_FPU.vhd:2877:57  */
  assign n4216 = n4199 & n4195;
  /* TG68K_FPU.vhd:2877:57  */
  assign n4217 = n4199 & n4195;
  /* TG68K_FPU.vhd:2788:57  */
  assign n4220 = n4079 ? n4186 : n4207;
  /* TG68K_FPU.vhd:2788:57  */
  assign n4221 = n4079 ? n4187 : n4208;
  /* TG68K_FPU.vhd:2788:57  */
  assign n4222 = n4079 ? n4188 : n4209;
  /* TG68K_FPU.vhd:2788:57  */
  assign n4223 = n4079 ? n4190 : n4211;
  /* TG68K_FPU.vhd:550:33  */
  assign n4230 = result_data[79]; // extract
  /* TG68K_FPU.vhd:551:37  */
  assign n4232 = result_data[78:64]; // extract
  /* TG68K_FPU.vhd:552:37  */
  assign n4234 = result_data[63:0]; // extract
  /* TG68K_FPU.vhd:558:29  */
  assign n4238 = n4232 == 15'b111111111111111;
  /* TG68K_FPU.vhd:560:36  */
  assign n4239 = result_data[63]; // extract
  /* TG68K_FPU.vhd:560:41  */
  assign n4240 = ~n4239;
  /* TG68K_FPU.vhd:560:58  */
  assign n4241 = result_data[62:0]; // extract
  /* TG68K_FPU.vhd:560:72  */
  assign n4243 = n4241 != 63'b000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:560:47  */
  assign n4244 = n4240 | n4243;
  assign n4247 = n4236[0]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n4248 = n4244 ? 1'b1 : n4247;
  assign n4249 = n4236[1]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n4250 = n4244 ? n4249 : 1'b1;
  assign n4251 = n4236[3]; // extract
  /* TG68K_FPU.vhd:560:25  */
  assign n4252 = n4244 ? n4251 : n4230;
  /* TG68K_FPU.vhd:568:32  */
  assign n4254 = n4232 == 15'b000000000000000;
  /* TG68K_FPU.vhd:568:68  */
  assign n4256 = n4234 == 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:568:55  */
  assign n4257 = n4256 & n4254;
  assign n4259 = {n4230, 1'b1};
  assign n4260 = n4259[0]; // extract
  assign n4261 = n4236[2]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n4262 = n4257 ? n4260 : n4261;
  assign n4263 = n4259[1]; // extract
  /* TG68K_FPU.vhd:568:17  */
  assign n4264 = n4257 ? n4263 : n4230;
  assign n4265 = {n4264, n4262};
  assign n4266 = {n4250, n4248};
  assign n4267 = n4236[1:0]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n4268 = n4238 ? n4266 : n4267;
  assign n4269 = n4265[0]; // extract
  assign n4270 = n4236[2]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n4271 = n4238 ? n4270 : n4269;
  assign n4272 = n4265[1]; // extract
  /* TG68K_FPU.vhd:558:17  */
  assign n4273 = n4238 ? n4252 : n4272;
  assign n4278 = fpsr[17]; // extract
  /* TG68K_FPU.vhd:2896:57  */
  assign n4279 = alu_overflow ? 1'b1 : n4278;
  assign n4280 = fpsr[25]; // extract
  /* TG68K_FPU.vhd:2896:57  */
  assign n4281 = alu_overflow ? 1'b1 : n4280;
  assign n4284 = fpsr[16]; // extract
  /* TG68K_FPU.vhd:2900:57  */
  assign n4285 = alu_underflow ? 1'b1 : n4284;
  assign n4286 = fpsr[24]; // extract
  /* TG68K_FPU.vhd:2900:57  */
  assign n4287 = alu_underflow ? 1'b1 : n4286;
  assign n4290 = fpsr[15]; // extract
  /* TG68K_FPU.vhd:2904:57  */
  assign n4291 = alu_inexact ? 1'b1 : n4290;
  assign n4292 = fpsr[23]; // extract
  /* TG68K_FPU.vhd:2904:57  */
  assign n4293 = alu_inexact ? 1'b1 : n4292;
  assign n4296 = fpsr[18]; // extract
  /* TG68K_FPU.vhd:2908:57  */
  assign n4297 = alu_invalid ? 1'b1 : n4296;
  assign n4298 = fpsr[26]; // extract
  /* TG68K_FPU.vhd:2908:57  */
  assign n4299 = alu_invalid ? 1'b1 : n4298;
  assign n4302 = fpsr[14]; // extract
  /* TG68K_FPU.vhd:2912:57  */
  assign n4303 = alu_divide_by_zero ? 1'b1 : n4302;
  assign n4304 = fpsr[22]; // extract
  /* TG68K_FPU.vhd:2912:57  */
  assign n4305 = alu_divide_by_zero ? 1'b1 : n4304;
  /* TG68K_FPU.vhd:2919:74  */
  assign n4307 = fpu_operation == 7'b0100001;
  /* TG68K_FPU.vhd:2919:101  */
  assign n4309 = fpu_operation == 7'b0100101;
  /* TG68K_FPU.vhd:2919:84  */
  assign n4310 = n4307 | n4309;
  /* TG68K_FPU.vhd:2922:98  */
  assign n4311 = result_data[6:0]; // extract
  assign n4312 = fpsr[21:19]; // extract
  assign n4313 = {n4293, n4305, n4312, n4297, n4279};
  /* TG68K_FPU.vhd:2919:57  */
  assign n4314 = n4310 ? n4311 : n4313;
  /* TG68K_FPU.vhd:2926:72  */
  assign n4316 = data_format == 3'b001;
  /* TG68K_FPU.vhd:2926:103  */
  assign n4318 = data_format == 3'b000;
  /* TG68K_FPU.vhd:2926:88  */
  assign n4319 = n4316 | n4318;
  /* TG68K_FPU.vhd:2927:92  */
  assign n4320 = result_data[31:0]; // extract
  /* TG68K_FPU.vhd:2928:75  */
  assign n4322 = data_format == 3'b101;
  /* TG68K_FPU.vhd:2929:92  */
  assign n4323 = result_data[63:32]; // extract
  /* TG68K_FPU.vhd:2928:57  */
  assign n4325 = n4322 ? n4323 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:2926:57  */
  assign n4326 = n4319 ? n4320 : n4325;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4327 = n4049 ? n6841 : n4326;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4329 = n4049 ? n4067 : 1'b1;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4330 = constrom_valid & n4049;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4333 = n4049 ? n4057 : n4220;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4334 = n4049 ? n4058 : n4221;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4335 = n4049 ? n4059 : n4222;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4336 = n4049 ? n4061 : n4223;
  assign n4337 = {n4299, n4281, n4287, n4314, n4285, n4291, n4303};
  assign n4338 = {n4273, n4271, n4268};
  assign n4339 = fpsr[26:14]; // extract
  /* TG68K_FPU.vhd:2766:49  */
  assign n4340 = n4049 ? n4339 : n4337;
  assign n4341 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:2766:49  */
  assign n4342 = n4049 ? n4341 : n4338;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4344 = n4049 ? n4074 : 4'b0000;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4345 = constrom_valid & n4049;
  /* TG68K_FPU.vhd:2766:49  */
  assign n4346 = constrom_valid & n4049;
  /* TG68K_FPU.vhd:2764:41  */
  assign n4348 = fpu_state == 4'b0110;
  /* TG68K_FPU.vhd:2937:41  */
  assign n4350 = fpu_state == 4'b0111;
  /* TG68K_FPU.vhd:2958:57  */
  assign n4353 = exception_code_internal == 8'b00000010;
  /* TG68K_FPU.vhd:2960:57  */
  assign n4357 = exception_code_internal == 8'b00000101;
  /* TG68K_FPU.vhd:2963:57  */
  assign n4361 = exception_code_internal == 8'b00001010;
  /* TG68K_FPU.vhd:2966:57  */
  assign n4365 = exception_code_internal == 8'b00001011;
  /* TG68K_FPU.vhd:2969:57  */
  assign n4369 = exception_code_internal == 8'b00001100;
  /* TG68K_FPU.vhd:2972:57  */
  assign n4373 = exception_code_internal == 8'b00001101;
  /* TG68K_FPU.vhd:2975:57  */
  assign n4377 = exception_code_internal == 8'b00001110;
  /* TG68K_FPU.vhd:2978:57  */
  assign n4381 = exception_code_internal == 8'b00001111;
  assign n4383 = {n4381, n4377, n4373, n4369, n4365, n4361, n4357, n4353};
  assign n4384 = fpsr[13]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4385 = n4384;
      8'b01000000: n4385 = n4384;
      8'b00100000: n4385 = n4384;
      8'b00010000: n4385 = n4384;
      8'b00001000: n4385 = 1'b1;
      8'b00000100: n4385 = n4384;
      8'b00000010: n4385 = n4384;
      8'b00000001: n4385 = n4384;
      default: n4385 = n4384;
    endcase
  assign n4386 = fpsr[14]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4387 = n4386;
      8'b01000000: n4387 = n4386;
      8'b00100000: n4387 = n4386;
      8'b00010000: n4387 = n4386;
      8'b00001000: n4387 = n4386;
      8'b00000100: n4387 = n4386;
      8'b00000010: n4387 = 1'b1;
      8'b00000001: n4387 = n4386;
      default: n4387 = n4386;
    endcase
  assign n4388 = fpsr[15]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4389 = 1'b1;
      8'b01000000: n4389 = n4388;
      8'b00100000: n4389 = n4388;
      8'b00010000: n4389 = n4388;
      8'b00001000: n4389 = n4388;
      8'b00000100: n4389 = n4388;
      8'b00000010: n4389 = n4388;
      8'b00000001: n4389 = n4388;
      default: n4389 = n4388;
    endcase
  assign n4390 = fpsr[16]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4391 = n4390;
      8'b01000000: n4391 = 1'b1;
      8'b00100000: n4391 = n4390;
      8'b00010000: n4391 = n4390;
      8'b00001000: n4391 = n4390;
      8'b00000100: n4391 = n4390;
      8'b00000010: n4391 = n4390;
      8'b00000001: n4391 = n4390;
      default: n4391 = n4390;
    endcase
  assign n4392 = fpsr[17]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4393 = n4392;
      8'b01000000: n4393 = n4392;
      8'b00100000: n4393 = 1'b1;
      8'b00010000: n4393 = n4392;
      8'b00001000: n4393 = n4392;
      8'b00000100: n4393 = n4392;
      8'b00000010: n4393 = n4392;
      8'b00000001: n4393 = n4392;
      default: n4393 = n4392;
    endcase
  assign n4394 = fpsr[18]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4395 = n4394;
      8'b01000000: n4395 = n4394;
      8'b00100000: n4395 = n4394;
      8'b00010000: n4395 = 1'b1;
      8'b00001000: n4395 = n4394;
      8'b00000100: n4395 = 1'b1;
      8'b00000010: n4395 = n4394;
      8'b00000001: n4395 = n4394;
      default: n4395 = n4394;
    endcase
  assign n4396 = fpsr[21]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4397 = n4396;
      8'b01000000: n4397 = n4396;
      8'b00100000: n4397 = n4396;
      8'b00010000: n4397 = n4396;
      8'b00001000: n4397 = 1'b1;
      8'b00000100: n4397 = n4396;
      8'b00000010: n4397 = n4396;
      8'b00000001: n4397 = 1'b1;
      default: n4397 = n4396;
    endcase
  assign n4398 = fpsr[22]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4399 = n4398;
      8'b01000000: n4399 = n4398;
      8'b00100000: n4399 = n4398;
      8'b00010000: n4399 = n4398;
      8'b00001000: n4399 = n4398;
      8'b00000100: n4399 = n4398;
      8'b00000010: n4399 = 1'b1;
      8'b00000001: n4399 = n4398;
      default: n4399 = n4398;
    endcase
  assign n4400 = fpsr[23]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4401 = 1'b1;
      8'b01000000: n4401 = n4400;
      8'b00100000: n4401 = n4400;
      8'b00010000: n4401 = n4400;
      8'b00001000: n4401 = n4400;
      8'b00000100: n4401 = n4400;
      8'b00000010: n4401 = n4400;
      8'b00000001: n4401 = n4400;
      default: n4401 = n4400;
    endcase
  assign n4402 = fpsr[24]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4403 = n4402;
      8'b01000000: n4403 = 1'b1;
      8'b00100000: n4403 = n4402;
      8'b00010000: n4403 = n4402;
      8'b00001000: n4403 = n4402;
      8'b00000100: n4403 = n4402;
      8'b00000010: n4403 = n4402;
      8'b00000001: n4403 = n4402;
      default: n4403 = n4402;
    endcase
  assign n4404 = fpsr[25]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4405 = n4404;
      8'b01000000: n4405 = n4404;
      8'b00100000: n4405 = 1'b1;
      8'b00010000: n4405 = n4404;
      8'b00001000: n4405 = n4404;
      8'b00000100: n4405 = n4404;
      8'b00000010: n4405 = n4404;
      8'b00000001: n4405 = n4404;
      default: n4405 = n4404;
    endcase
  assign n4406 = fpsr[26]; // extract
  /* TG68K_FPU.vhd:2957:49  */
  always @*
    case (n4383)
      8'b10000000: n4407 = n4406;
      8'b01000000: n4407 = n4406;
      8'b00100000: n4407 = n4406;
      8'b00010000: n4407 = 1'b1;
      8'b00001000: n4407 = n4406;
      8'b00000100: n4407 = 1'b1;
      8'b00000010: n4407 = n4406;
      8'b00000001: n4407 = n4406;
      default: n4407 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:2989:72  */
  assign n4408 = fpcr[15]; // extract
  /* TG68K_FPU.vhd:2989:65  */
  assign n4411 = n4408 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:2988:57  */
  assign n4413 = exception_code_internal == 8'b00000010;
  /* TG68K_FPU.vhd:2995:72  */
  assign n4414 = fpcr[10]; // extract
  /* TG68K_FPU.vhd:2995:65  */
  assign n4417 = n4414 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:2994:57  */
  assign n4419 = exception_code_internal == 8'b00000101;
  /* TG68K_FPU.vhd:3001:72  */
  assign n4420 = fpcr[13]; // extract
  /* TG68K_FPU.vhd:3001:65  */
  assign n4423 = n4420 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:3000:57  */
  assign n4425 = exception_code_internal == 8'b00001100;
  /* TG68K_FPU.vhd:3007:72  */
  assign n4426 = fpcr[12]; // extract
  /* TG68K_FPU.vhd:3007:65  */
  assign n4429 = n4426 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:3006:57  */
  assign n4431 = exception_code_internal == 8'b00001101;
  /* TG68K_FPU.vhd:3013:72  */
  assign n4432 = fpcr[11]; // extract
  /* TG68K_FPU.vhd:3013:65  */
  assign n4435 = n4432 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:3012:57  */
  assign n4437 = exception_code_internal == 8'b00001110;
  /* TG68K_FPU.vhd:3019:72  */
  assign n4438 = fpcr[9]; // extract
  /* TG68K_FPU.vhd:3019:65  */
  assign n4441 = n4438 ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:3018:57  */
  assign n4443 = exception_code_internal == 8'b00001111;
  assign n4444 = {n4443, n4437, n4431, n4425, n4419, n4413};
  /* TG68K_FPU.vhd:2987:49  */
  always @*
    case (n4444)
      6'b100000: n4446 = n4441;
      6'b010000: n4446 = n4435;
      6'b001000: n4446 = n4429;
      6'b000100: n4446 = n4423;
      6'b000010: n4446 = n4417;
      6'b000001: n4446 = n4411;
      default: n4446 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:2947:41  */
  assign n4448 = fpu_state == 4'b1000;
  /* TG68K_FPU.vhd:3044:116  */
  assign n4450 = {fsave_frame_format_latched, 24'b000000000000000000000000};
  /* TG68K_FPU.vhd:3040:65  */
  assign n4452 = fsave_data_index == 6'b000000;
  /* TG68K_FPU.vhd:3047:103  */
  assign n4454 = fsave_frame_format_latched == 8'b00000000;
  /* TG68K_FPU.vhd:3047:73  */
  assign n4456 = n4454 ? 32'b00000000000000000000000000000000 : fpiar;
  /* TG68K_FPU.vhd:3045:65  */
  assign n4458 = fsave_data_index == 6'b000001;
  /* TG68K_FPU.vhd:3056:103  */
  assign n4460 = fsave_frame_format_latched == 8'b01100000;
  /* TG68K_FPU.vhd:3056:141  */
  assign n4462 = fsave_frame_format_latched == 8'b11011000;
  /* TG68K_FPU.vhd:3056:111  */
  assign n4463 = n4460 | n4462;
  /* TG68K_FPU.vhd:3056:73  */
  assign n4465 = n4463 ? fpcr : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:3054:65  */
  assign n4467 = fsave_data_index == 6'b000010;
  /* TG68K_FPU.vhd:3063:103  */
  assign n4469 = fsave_frame_format_latched == 8'b01100000;
  /* TG68K_FPU.vhd:3063:141  */
  assign n4471 = fsave_frame_format_latched == 8'b11011000;
  /* TG68K_FPU.vhd:3063:111  */
  assign n4472 = n4469 | n4471;
  /* TG68K_FPU.vhd:3063:73  */
  assign n4474 = n4472 ? fpsr : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:3061:65  */
  assign n4476 = fsave_data_index == 6'b000011;
  /* TG68K_FPU.vhd:3068:65  */
  assign n4479 = $unsigned(fsave_data_index) >= $unsigned(6'b000100);
  /* TG68K_FPU.vhd:3068:65  */
  assign n4480 = $unsigned(fsave_data_index) <= $unsigned(6'b011011);
  /* TG68K_FPU.vhd:3068:65  */
  assign n4481 = n4479 & n4480;
  /* TG68K_FPU.vhd:3074:103  */
  assign n4483 = fsave_frame_format_latched == 8'b11011000;
  /* TG68K_FPU.vhd:3075:127  */
  assign n4484 = {26'b0, fsave_data_index};  //  uext
  /* TG68K_FPU.vhd:3075:127  */
  assign n4486 = n4484 - 32'b00000000000000000000000000011100;
  /* TG68K_FPU.vhd:3075:127  */
  assign n4487 = n4486[2:0];  // trunc
  /* TG68K_FPU.vhd:3075:127  */
  assign n4489 = 3'b111 - n4487;
  /* TG68K_FPU.vhd:3075:132  */
  assign n4491 = fp_registers[n6963 + 48 +: 32]; //(dyn_extract)
  /* TG68K_FPU.vhd:3074:73  */
  assign n4493 = n4483 ? n4491 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:3072:65  */
  assign n4496 = $unsigned(fsave_data_index) >= $unsigned(6'b011100);
  /* TG68K_FPU.vhd:3072:65  */
  assign n4497 = $unsigned(fsave_data_index) <= $unsigned(6'b100011);
  /* TG68K_FPU.vhd:3072:65  */
  assign n4498 = n4496 & n4497;
  /* TG68K_FPU.vhd:3081:103  */
  assign n4500 = fsave_frame_format_latched == 8'b11011000;
  /* TG68K_FPU.vhd:3082:127  */
  assign n4501 = {26'b0, fsave_data_index};  //  uext
  /* TG68K_FPU.vhd:3082:127  */
  assign n4503 = n4501 - 32'b00000000000000000000000000100100;
  /* TG68K_FPU.vhd:3082:127  */
  assign n4504 = n4503[2:0];  // trunc
  /* TG68K_FPU.vhd:3082:127  */
  assign n4506 = 3'b111 - n4504;
  /* TG68K_FPU.vhd:3082:132  */
  assign n4508 = fp_registers[n6966 + 16 +: 32]; //(dyn_extract)
  /* TG68K_FPU.vhd:3081:73  */
  assign n4510 = n4500 ? n4508 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:3079:65  */
  assign n4513 = $unsigned(fsave_data_index) >= $unsigned(6'b100100);
  /* TG68K_FPU.vhd:3079:65  */
  assign n4514 = $unsigned(fsave_data_index) <= $unsigned(6'b101011);
  /* TG68K_FPU.vhd:3079:65  */
  assign n4515 = n4513 & n4514;
  /* TG68K_FPU.vhd:3089:103  */
  assign n4517 = fsave_frame_format_latched == 8'b11011000;
  /* TG68K_FPU.vhd:3090:141  */
  assign n4518 = {26'b0, fsave_data_index};  //  uext
  /* TG68K_FPU.vhd:3090:141  */
  assign n4520 = n4518 - 32'b00000000000000000000000000101100;
  /* TG68K_FPU.vhd:3090:141  */
  assign n4521 = n4520[2:0];  // trunc
  /* TG68K_FPU.vhd:3090:141  */
  assign n4523 = 3'b111 - n4521;
  assign n4527 = {n6968, 16'b0000000000000000};
  /* TG68K_FPU.vhd:3089:73  */
  assign n4529 = n4517 ? n4527 : 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:3086:65  */
  assign n4532 = $unsigned(fsave_data_index) >= $unsigned(6'b101100);
  /* TG68K_FPU.vhd:3086:65  */
  assign n4533 = $unsigned(fsave_data_index) <= $unsigned(6'b110011);
  /* TG68K_FPU.vhd:3086:65  */
  assign n4534 = n4532 & n4533;
  /* TG68K_FPU.vhd:3095:65  */
  assign n4539 = $unsigned(fsave_data_index) >= $unsigned(6'b110100);
  /* TG68K_FPU.vhd:3095:65  */
  assign n4540 = $unsigned(fsave_data_index) <= $unsigned(6'b110101);
  /* TG68K_FPU.vhd:3095:65  */
  assign n4541 = n4539 & n4540;
  assign n4542 = {n4541, n4534, n4515, n4498, n4481, n4476, n4467, n4458, n4452};
  /* TG68K_FPU.vhd:3039:57  */
  always @*
    case (n4542)
      9'b100000000: n4546 = 32'b00000000000000000000000000000000;
      9'b010000000: n4546 = n4529;
      9'b001000000: n4546 = n4510;
      9'b000100000: n4546 = n4493;
      9'b000010000: n4546 = 32'b00000000000000000000000000000000;
      9'b000001000: n4546 = n4474;
      9'b000000100: n4546 = n4465;
      9'b000000010: n4546 = n4456;
      9'b000000001: n4546 = n4450;
      default: n4546 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:3038:49  */
  assign n4547 = fsave_data_request ? n4546 : n6841;
  /* TG68K_FPU.vhd:3112:114  */
  assign n4548 = {26'b0, fsave_data_index};  //  uext
  /* TG68K_FPU.vhd:3112:114  */
  assign n4550 = n4548 == 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:3112:93  */
  assign n4551 = n4550 & fsave_data_request;
  /* TG68K_FPU.vhd:3112:65  */
  assign n4553 = n4551 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3112:65  */
  assign n4555 = n4551 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3110:57  */
  assign n4557 = fsave_frame_format_latched == 8'b00000000;
  /* TG68K_FPU.vhd:3119:114  */
  assign n4558 = {26'b0, fsave_data_index};  //  uext
  /* TG68K_FPU.vhd:3119:114  */
  assign n4560 = n4558 == 32'b00000000000000000000000000001110;
  /* TG68K_FPU.vhd:3119:93  */
  assign n4561 = n4560 & fsave_data_request;
  /* TG68K_FPU.vhd:3119:65  */
  assign n4563 = n4561 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3119:65  */
  assign n4565 = n4561 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3117:57  */
  assign n4567 = fsave_frame_format_latched == 8'b01100000;
  /* TG68K_FPU.vhd:3126:114  */
  assign n4568 = {26'b0, fsave_data_index};  //  uext
  /* TG68K_FPU.vhd:3126:114  */
  assign n4570 = n4568 == 32'b00000000000000000000000000110101;
  /* TG68K_FPU.vhd:3126:93  */
  assign n4571 = n4570 & fsave_data_request;
  /* TG68K_FPU.vhd:3126:65  */
  assign n4573 = n4571 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3126:65  */
  assign n4575 = n4571 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3124:57  */
  assign n4577 = fsave_frame_format_latched == 8'b11011000;
  /* TG68K_FPU.vhd:3133:114  */
  assign n4578 = {26'b0, fsave_data_index};  //  uext
  /* TG68K_FPU.vhd:3133:114  */
  assign n4580 = n4578 == 32'b00000000000000000000000000001110;
  /* TG68K_FPU.vhd:3133:93  */
  assign n4581 = n4580 & fsave_data_request;
  /* TG68K_FPU.vhd:3133:65  */
  assign n4583 = n4581 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3133:65  */
  assign n4585 = n4581 ? 4'b0000 : fpu_state;
  assign n4586 = {n4577, n4567, n4557};
  /* TG68K_FPU.vhd:3109:49  */
  always @*
    case (n4586)
      3'b100: n4587 = n4573;
      3'b010: n4587 = n4563;
      3'b001: n4587 = n4553;
      default: n4587 = n4583;
    endcase
  /* TG68K_FPU.vhd:3109:49  */
  always @*
    case (n4586)
      3'b100: n4588 = n4575;
      3'b010: n4588 = n4565;
      3'b001: n4588 = n4555;
      default: n4588 = n4585;
    endcase
  /* TG68K_FPU.vhd:3034:41  */
  assign n4590 = fpu_state == 4'b1001;
  /* TG68K_FPU.vhd:3150:114  */
  assign n4591 = frestore_data_in[31:24]; // extract
  /* TG68K_FPU.vhd:3151:94  */
  assign n4592 = frestore_data_in[31:24]; // extract
  /* TG68K_FPU.vhd:3152:81  */
  assign n4602 = n4592 == 8'b00000000;
  /* TG68K_FPU.vhd:3168:81  */
  assign n4604 = n4592 == 8'b00000001;
  /* TG68K_FPU.vhd:3176:120  */
  assign n4605 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3176:120  */
  assign n4607 = n4605 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3176:106  */
  assign n4608 = n4607[5:0];  // trunc
  /* TG68K_FPU.vhd:3174:81  */
  assign n4610 = n4592 == 8'b00011000;
  /* TG68K_FPU.vhd:3180:120  */
  assign n4611 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3180:120  */
  assign n4613 = n4611 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3180:106  */
  assign n4614 = n4613[5:0];  // trunc
  /* TG68K_FPU.vhd:3178:81  */
  assign n4616 = n4592 == 8'b01000001;
  /* TG68K_FPU.vhd:3184:120  */
  assign n4617 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3184:120  */
  assign n4619 = n4617 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3184:106  */
  assign n4620 = n4619[5:0];  // trunc
  /* TG68K_FPU.vhd:3182:81  */
  assign n4622 = n4592 == 8'b01100000;
  /* TG68K_FPU.vhd:3188:120  */
  assign n4623 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3188:120  */
  assign n4625 = n4623 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3188:106  */
  assign n4626 = n4625[5:0];  // trunc
  /* TG68K_FPU.vhd:3186:81  */
  assign n4628 = n4592 == 8'b00111000;
  assign n4629 = {n4628, n4622, n4616, n4610, n4604, n4602};
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4632 = fpu_done_i;
      6'b010000: n4632 = fpu_done_i;
      6'b001000: n4632 = fpu_done_i;
      6'b000100: n4632 = fpu_done_i;
      6'b000010: n4632 = 1'b1;
      6'b000001: n4632 = 1'b1;
      default: n4632 = fpu_done_i;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4634 = fpu_exception_i;
      6'b010000: n4634 = fpu_exception_i;
      6'b001000: n4634 = fpu_exception_i;
      6'b000100: n4634 = fpu_exception_i;
      6'b000010: n4634 = fpu_exception_i;
      6'b000001: n4634 = fpu_exception_i;
      default: n4634 = 1'b1;
    endcase
  assign n4635 = n755[79:0]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4636 = n4635;
      6'b010000: n4636 = n4635;
      6'b001000: n4636 = n4635;
      6'b000100: n4636 = n4635;
      6'b000010: n4636 = n4635;
      6'b000001: n4636 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4636 = n4635;
    endcase
  assign n4637 = n755[159:80]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4638 = n4637;
      6'b010000: n4638 = n4637;
      6'b001000: n4638 = n4637;
      6'b000100: n4638 = n4637;
      6'b000010: n4638 = n4637;
      6'b000001: n4638 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4638 = n4637;
    endcase
  assign n4639 = n755[239:160]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4640 = n4639;
      6'b010000: n4640 = n4639;
      6'b001000: n4640 = n4639;
      6'b000100: n4640 = n4639;
      6'b000010: n4640 = n4639;
      6'b000001: n4640 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4640 = n4639;
    endcase
  assign n4641 = n755[319:240]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4642 = n4641;
      6'b010000: n4642 = n4641;
      6'b001000: n4642 = n4641;
      6'b000100: n4642 = n4641;
      6'b000010: n4642 = n4641;
      6'b000001: n4642 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4642 = n4641;
    endcase
  assign n4643 = n755[399:320]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4644 = n4643;
      6'b010000: n4644 = n4643;
      6'b001000: n4644 = n4643;
      6'b000100: n4644 = n4643;
      6'b000010: n4644 = n4643;
      6'b000001: n4644 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4644 = n4643;
    endcase
  assign n4645 = n755[479:400]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4646 = n4645;
      6'b010000: n4646 = n4645;
      6'b001000: n4646 = n4645;
      6'b000100: n4646 = n4645;
      6'b000010: n4646 = n4645;
      6'b000001: n4646 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4646 = n4645;
    endcase
  assign n4647 = n755[559:480]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4648 = n4647;
      6'b010000: n4648 = n4647;
      6'b001000: n4648 = n4647;
      6'b000100: n4648 = n4647;
      6'b000010: n4648 = n4647;
      6'b000001: n4648 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4648 = n4647;
    endcase
  assign n4649 = n755[639:560]; // extract
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4650 = n4649;
      6'b010000: n4650 = n4649;
      6'b001000: n4650 = n4649;
      6'b000100: n4650 = n4649;
      6'b000010: n4650 = n4649;
      6'b000001: n4650 = 80'b01111111111111111100000000000000000000000000000000000000000000000000000000000000;
      default: n4650 = n4649;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4652 = fpcr;
      6'b010000: n4652 = fpcr;
      6'b001000: n4652 = fpcr;
      6'b000100: n4652 = fpcr;
      6'b000010: n4652 = fpcr;
      6'b000001: n4652 = 32'b00000000000000000000000000000000;
      default: n4652 = fpcr;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4654 = fpsr;
      6'b010000: n4654 = fpsr;
      6'b001000: n4654 = fpsr;
      6'b000100: n4654 = fpsr;
      6'b000010: n4654 = fpsr;
      6'b000001: n4654 = 32'b00000000000000000000000000000000;
      default: n4654 = fpsr;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4656 = fpiar;
      6'b010000: n4656 = fpiar;
      6'b001000: n4656 = fpiar;
      6'b000100: n4656 = fpiar;
      6'b000010: n4656 = fpiar;
      6'b000001: n4656 = 32'b00000000000000000000000000000000;
      default: n4656 = fpiar;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4660 = fpu_state;
      6'b010000: n4660 = fpu_state;
      6'b001000: n4660 = fpu_state;
      6'b000100: n4660 = fpu_state;
      6'b000010: n4660 = 4'b0000;
      6'b000001: n4660 = 4'b0000;
      default: n4660 = 4'b1000;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4662 = fpu_just_reset;
      6'b010000: n4662 = fpu_just_reset;
      6'b001000: n4662 = fpu_just_reset;
      6'b000100: n4662 = fpu_just_reset;
      6'b000010: n4662 = fpu_just_reset;
      6'b000001: n4662 = 1'b1;
      default: n4662 = fpu_just_reset;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4663 = n4626;
      6'b010000: n4663 = n4620;
      6'b001000: n4663 = n4614;
      6'b000100: n4663 = n4608;
      6'b000010: n4663 = fsave_counter;
      6'b000001: n4663 = fsave_counter;
      default: n4663 = fsave_counter;
    endcase
  /* TG68K_FPU.vhd:3151:73  */
  always @*
    case (n4629)
      6'b100000: n4665 = exception_code_internal;
      6'b010000: n4665 = exception_code_internal;
      6'b001000: n4665 = exception_code_internal;
      6'b000100: n4665 = exception_code_internal;
      6'b000010: n4665 = exception_code_internal;
      6'b000001: n4665 = exception_code_internal;
      default: n4665 = 8'b00001010;
    endcase
  /* TG68K_FPU.vhd:3148:65  */
  assign n4667 = fsave_counter == 6'b000000;
  /* TG68K_FPU.vhd:3200:104  */
  assign n4668 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3200:104  */
  assign n4670 = n4668 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3200:90  */
  assign n4671 = n4670[5:0];  // trunc
  /* TG68K_FPU.vhd:3197:65  */
  assign n4673 = fsave_counter == 6'b000001;
  /* TG68K_FPU.vhd:613:28  */
  assign n4679 = frestore_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:613:41  */
  assign n4681 = n4679 == 2'b11;
  /* TG68K_FPU.vhd:613:17  */
  assign n4685 = n4681 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:613:17  */
  assign n4691 = n4681 ? 1'b0 : 1'bX;
  /* TG68K_FPU.vhd:618:28  */
  assign n4692 = frestore_data_in[31:16]; // extract
  /* TG68K_FPU.vhd:618:43  */
  assign n4694 = n4692 != 16'b0000000000000000;
  /* TG68K_FPU.vhd:618:65  */
  assign n4695 = frestore_data_in[5:0]; // extract
  /* TG68K_FPU.vhd:618:78  */
  assign n4697 = n4695 != 6'b000000;
  /* TG68K_FPU.vhd:618:54  */
  assign n4698 = n4694 | n4697;
  /* TG68K_FPU.vhd:618:17  */
  assign n4701 = n4708 ? 1'b0 : n4685;
  /* TG68K_FPU.vhd:618:17  */
  assign n4704 = n4710 ? 1'b0 : n4691;
  /* TG68K_FPU.vhd:618:17  */
  assign n4705 = n4685 & n4698;
  /* TG68K_FPU.vhd:618:17  */
  assign n4707 = n4685 & n4698;
  /* TG68K_FPU.vhd:618:17  */
  assign n4708 = n4705 & n4685;
  /* TG68K_FPU.vhd:618:17  */
  assign n4710 = n4707 & n4685;
  /* TG68K_FPU.vhd:623:17  */
  assign n4716 = n4701 ? 1'b1 : n4704;
  /* TG68K_FPU.vhd:597:30  */
  assign n4724 = frestore_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:43  */
  assign n4726 = n4724 == 2'b11;
  assign n4728 = frestore_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:17  */
  assign n4729 = n4726 ? 2'b00 : n4728;
  assign n4733 = frestore_data_in[15:8]; // extract
  assign n4735 = {16'b0000000000000000, n4733, n4729, 6'b000000};
  /* TG68K_FPU.vhd:597:30  */
  assign n4743 = frestore_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:43  */
  assign n4745 = n4743 == 2'b11;
  assign n4747 = frestore_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:17  */
  assign n4748 = n4745 ? 2'b00 : n4747;
  assign n4752 = frestore_data_in[15:8]; // extract
  assign n4754 = {16'b0000000000000000, n4752, n4748, 6'b000000};
  /* TG68K_FPU.vhd:3213:100  */
  assign n4755 = frestore_data_in[15:14]; // extract
  /* TG68K_FPU.vhd:3213:115  */
  assign n4757 = n4755 == 2'b11;
  /* TG68K_FPU.vhd:3213:81  */
  assign n4760 = n4757 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:3218:100  */
  assign n4761 = frestore_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:3218:113  */
  assign n4763 = n4761 == 2'b11;
  /* TG68K_FPU.vhd:3218:81  */
  assign n4766 = n4763 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:3204:73  */
  assign n4767 = n4716 ? n4735 : n4754;
  /* TG68K_FPU.vhd:3204:73  */
  assign n4772 = n4716 ? 1'b1 : n4760;
  /* TG68K_FPU.vhd:3204:73  */
  assign n4774 = n4716 ? 1'b1 : n4766;
  /* TG68K_FPU.vhd:3224:104  */
  assign n4775 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3224:104  */
  assign n4777 = n4775 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3224:90  */
  assign n4778 = n4777[5:0];  // trunc
  /* TG68K_FPU.vhd:3202:65  */
  assign n4780 = fsave_counter == 6'b000010;
  /* TG68K_FPU.vhd:3233:81  */
  assign n4789 = frestore_frame_format == 8'b00011000;
  /* TG68K_FPU.vhd:3240:120  */
  assign n4790 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3240:120  */
  assign n4792 = n4790 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3240:106  */
  assign n4793 = n4792[5:0];  // trunc
  /* TG68K_FPU.vhd:3237:81  */
  assign n4795 = frestore_frame_format == 8'b01000001;
  /* TG68K_FPU.vhd:3237:92  */
  assign n4797 = frestore_frame_format == 8'b01100000;
  /* TG68K_FPU.vhd:3237:92  */
  assign n4798 = n4795 | n4797;
  /* TG68K_FPU.vhd:3243:120  */
  assign n4799 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3243:120  */
  assign n4801 = n4799 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3243:106  */
  assign n4802 = n4801[5:0];  // trunc
  /* TG68K_FPU.vhd:3241:81  */
  assign n4804 = frestore_frame_format == 8'b00111000;
  /* TG68K_FPU.vhd:3246:120  */
  assign n4805 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3246:120  */
  assign n4807 = n4805 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3246:106  */
  assign n4808 = n4807[5:0];  // trunc
  /* TG68K_FPU.vhd:3244:81  */
  assign n4810 = frestore_frame_format == 8'b11011000;
  assign n4811 = {n4810, n4804, n4798, n4789};
  /* TG68K_FPU.vhd:3232:73  */
  always @*
    case (n4811)
      4'b1000: n4814 = fpu_done_i;
      4'b0100: n4814 = fpu_done_i;
      4'b0010: n4814 = fpu_done_i;
      4'b0001: n4814 = 1'b1;
      default: n4814 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:3232:73  */
  always @*
    case (n4811)
      4'b1000: n4817 = fpu_state;
      4'b0100: n4817 = fpu_state;
      4'b0010: n4817 = fpu_state;
      4'b0001: n4817 = 4'b0000;
      default: n4817 = 4'b0000;
    endcase
  /* TG68K_FPU.vhd:3232:73  */
  always @*
    case (n4811)
      4'b1000: n4818 = n4808;
      4'b0100: n4818 = n4802;
      4'b0010: n4818 = n4793;
      4'b0001: n4818 = fsave_counter;
      default: n4818 = fsave_counter;
    endcase
  /* TG68K_FPU.vhd:3226:65  */
  assign n4820 = fsave_counter == 6'b000011;
  /* TG68K_FPU.vhd:3257:98  */
  assign n4822 = frestore_frame_format == 8'b01000001;
  /* TG68K_FPU.vhd:3257:131  */
  assign n4824 = frestore_frame_format == 8'b01100000;
  /* TG68K_FPU.vhd:3257:106  */
  assign n4825 = n4822 | n4824;
  /* TG68K_FPU.vhd:3258:98  */
  assign n4826 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3258:98  */
  assign n4828 = n4826 == 32'b00000000000000000000000000001110;
  /* TG68K_FPU.vhd:3263:120  */
  assign n4829 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3263:120  */
  assign n4831 = n4829 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3263:106  */
  assign n4832 = n4831[5:0];  // trunc
  /* TG68K_FPU.vhd:3257:73  */
  assign n4834 = n4842 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3257:73  */
  assign n4836 = n4843 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3258:81  */
  assign n4837 = n4828 ? fsave_counter : n4832;
  /* TG68K_FPU.vhd:3267:112  */
  assign n4838 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3267:112  */
  assign n4840 = n4838 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3267:98  */
  assign n4841 = n4840[5:0];  // trunc
  /* TG68K_FPU.vhd:3257:73  */
  assign n4842 = n4828 & n4825;
  /* TG68K_FPU.vhd:3257:73  */
  assign n4843 = n4828 & n4825;
  /* TG68K_FPU.vhd:3257:73  */
  assign n4844 = n4825 ? n4837 : n4841;
  /* TG68K_FPU.vhd:3253:65  */
  assign n4847 = $unsigned(fsave_counter) >= $unsigned(6'b000100);
  /* TG68K_FPU.vhd:3253:65  */
  assign n4848 = $unsigned(fsave_counter) <= $unsigned(6'b001110);
  /* TG68K_FPU.vhd:3253:65  */
  assign n4849 = n4847 & n4848;
  /* TG68K_FPU.vhd:3273:104  */
  assign n4850 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3273:104  */
  assign n4852 = n4850 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3273:90  */
  assign n4853 = n4852[5:0];  // trunc
  /* TG68K_FPU.vhd:3270:65  */
  assign n4856 = $unsigned(fsave_counter) >= $unsigned(6'b001111);
  /* TG68K_FPU.vhd:3270:65  */
  assign n4857 = $unsigned(fsave_counter) <= $unsigned(6'b011011);
  /* TG68K_FPU.vhd:3270:65  */
  assign n4858 = n4856 & n4857;
  /* TG68K_FPU.vhd:3280:106  */
  assign n4859 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3280:106  */
  assign n4861 = n4859 == 32'b00000000000000000000000000010111;
  /* TG68K_FPU.vhd:3285:128  */
  assign n4862 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3285:128  */
  assign n4864 = n4862 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3285:114  */
  assign n4865 = n4864[5:0];  // trunc
  /* TG68K_FPU.vhd:3280:89  */
  assign n4867 = n4861 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3280:89  */
  assign n4869 = n4861 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3280:89  */
  assign n4870 = n4861 ? fsave_counter : n4865;
  /* TG68K_FPU.vhd:3278:81  */
  assign n4872 = frestore_frame_format == 8'b00111000;
  /* TG68K_FPU.vhd:3295:136  */
  assign n4873 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3295:136  */
  assign n4875 = n4873 - 32'b00000000000000000000000000011100;
  /* TG68K_FPU.vhd:3295:136  */
  assign n4876 = n4875[2:0];  // trunc
  /* TG68K_FPU.vhd:3295:136  */
  assign n4878 = 3'b111 - n4876;
  /* TG68K_FPU.vhd:3296:136  */
  assign n4881 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3296:136  */
  assign n4883 = n4881 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3296:122  */
  assign n4884 = n4883[5:0];  // trunc
  /* TG68K_FPU.vhd:3291:97  */
  assign n4887 = $unsigned(fsave_counter) >= $unsigned(6'b011100);
  /* TG68K_FPU.vhd:3291:97  */
  assign n4888 = $unsigned(fsave_counter) <= $unsigned(6'b100011);
  /* TG68K_FPU.vhd:3291:97  */
  assign n4889 = n4887 & n4888;
  /* TG68K_FPU.vhd:3301:136  */
  assign n4890 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3301:136  */
  assign n4892 = n4890 - 32'b00000000000000000000000000100100;
  /* TG68K_FPU.vhd:3301:136  */
  assign n4893 = n4892[2:0];  // trunc
  /* TG68K_FPU.vhd:3301:136  */
  assign n4895 = 3'b111 - n4893;
  /* TG68K_FPU.vhd:3302:136  */
  assign n4898 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3302:136  */
  assign n4900 = n4898 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3302:122  */
  assign n4901 = n4900[5:0];  // trunc
  /* TG68K_FPU.vhd:3297:97  */
  assign n4904 = $unsigned(fsave_counter) >= $unsigned(6'b100100);
  /* TG68K_FPU.vhd:3297:97  */
  assign n4905 = $unsigned(fsave_counter) <= $unsigned(6'b101011);
  /* TG68K_FPU.vhd:3297:97  */
  assign n4906 = n4904 & n4905;
  /* TG68K_FPU.vhd:3307:136  */
  assign n4907 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3307:136  */
  assign n4909 = n4907 - 32'b00000000000000000000000000101100;
  /* TG68K_FPU.vhd:3307:136  */
  assign n4910 = n4909[2:0];  // trunc
  /* TG68K_FPU.vhd:3307:136  */
  assign n4912 = 3'b111 - n4910;
  /* TG68K_FPU.vhd:3307:174  */
  assign n4914 = frestore_data_in[31:16]; // extract
  /* TG68K_FPU.vhd:3309:169  */
  assign n4916 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3309:169  */
  assign n4918 = n4916 - 32'b00000000000000000000000000101100;
  /* TG68K_FPU.vhd:3309:155  */
  assign n4919 = n4918[30:0];  // trunc
  /* TG68K_FPU.vhd:3309:143  */
  assign n4920 = n4919[2:0];  // trunc
  /* TG68K_FPU.vhd:3310:157  */
  assign n4921 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3310:157  */
  assign n4923 = n4921 - 32'b00000000000000000000000000101100;
  /* TG68K_FPU.vhd:3310:157  */
  assign n4924 = n4923[2:0];  // trunc
  /* TG68K_FPU.vhd:3310:157  */
  assign n4926 = 3'b111 - n4924;
  /* TG68K_FPU.vhd:3310:162  */
  assign n4928 = frestore_fp_temp[n7101 + 16 +: 64]; //(dyn_extract)
  /* TG68K_FPU.vhd:3310:195  */
  assign n4929 = frestore_data_in[31:16]; // extract
  /* TG68K_FPU.vhd:3310:177  */
  assign n4930 = {n4928, n4929};
  /* TG68K_FPU.vhd:3316:136  */
  assign n4943 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3316:136  */
  assign n4945 = n4943 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3316:122  */
  assign n4946 = n4945[5:0];  // trunc
  /* TG68K_FPU.vhd:3303:97  */
  assign n4949 = $unsigned(fsave_counter) >= $unsigned(6'b101100);
  /* TG68K_FPU.vhd:3303:97  */
  assign n4950 = $unsigned(fsave_counter) <= $unsigned(6'b110011);
  /* TG68K_FPU.vhd:3303:97  */
  assign n4951 = n4949 & n4950;
  /* TG68K_FPU.vhd:3320:122  */
  assign n4952 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3320:122  */
  assign n4954 = n4952 == 32'b00000000000000000000000000110101;
  /* TG68K_FPU.vhd:3325:144  */
  assign n4955 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3325:144  */
  assign n4957 = n4955 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3325:130  */
  assign n4958 = n4957[5:0];  // trunc
  /* TG68K_FPU.vhd:3320:105  */
  assign n4960 = n4954 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3320:105  */
  assign n4962 = n4954 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3320:105  */
  assign n4963 = n4954 ? fsave_counter : n4958;
  assign n4964 = {n4951, n4906, n4889};
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4965 = fpu_done_i;
      3'b010: n4965 = fpu_done_i;
      3'b001: n4965 = fpu_done_i;
      default: n4965 = n4960;
    endcase
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4970 = 1'b1;
      3'b010: n4970 = 1'b0;
      3'b001: n4970 = 1'b0;
      default: n4970 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4971 = n4920;
      3'b010: n4971 = fp_reg_write_addr;
      3'b001: n4971 = fp_reg_write_addr;
      default: n4971 = fp_reg_write_addr;
    endcase
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4972 = n4930;
      3'b010: n4972 = fp_reg_write_data;
      3'b001: n4972 = fp_reg_write_data;
      default: n4972 = fp_reg_write_data;
    endcase
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4975 = 1'b1;
      3'b010: n4975 = 1'b0;
      3'b001: n4975 = 1'b0;
      default: n4975 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4976 = fpu_state;
      3'b010: n4976 = fpu_state;
      3'b001: n4976 = fpu_state;
      default: n4976 = n4962;
    endcase
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4977 = n4946;
      3'b010: n4977 = n4901;
      3'b001: n4977 = n4884;
      default: n4977 = n4963;
    endcase
  /* TG68K_FPU.vhd:3290:89  */
  always @*
    case (n4964)
      3'b100: n4978 = n7098;
      3'b010: n4978 = n7055;
      3'b001: n4978 = n7011;
      default: n4978 = frestore_fp_temp;
    endcase
  /* TG68K_FPU.vhd:3287:81  */
  assign n4980 = frestore_frame_format == 8'b11011000;
  /* TG68K_FPU.vhd:3331:106  */
  assign n4981 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3331:106  */
  assign n4983 = n4981 == 32'b00000000000000000000000000110101;
  /* TG68K_FPU.vhd:3335:128  */
  assign n4984 = {26'b0, fsave_counter};  //  uext
  /* TG68K_FPU.vhd:3335:128  */
  assign n4986 = n4984 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3335:114  */
  assign n4987 = n4986[5:0];  // trunc
  /* TG68K_FPU.vhd:3331:89  */
  assign n4989 = n4983 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3331:89  */
  assign n4991 = n4983 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3331:89  */
  assign n4992 = n4983 ? fsave_counter : n4987;
  assign n4993 = {n4980, n4872};
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n4994 = n4965;
      2'b01: n4994 = n4867;
      default: n4994 = n4989;
    endcase
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n4998 = n4970;
      2'b01: n4998 = 1'b0;
      default: n4998 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n4999 = n4971;
      2'b01: n4999 = fp_reg_write_addr;
      default: n4999 = fp_reg_write_addr;
    endcase
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n5000 = n4972;
      2'b01: n5000 = fp_reg_write_data;
      default: n5000 = fp_reg_write_data;
    endcase
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n5002 = n4975;
      2'b01: n5002 = 1'b0;
      default: n5002 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n5003 = n4976;
      2'b01: n5003 = n4869;
      default: n5003 = n4991;
    endcase
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n5004 = n4977;
      2'b01: n5004 = n4870;
      default: n5004 = n4992;
    endcase
  /* TG68K_FPU.vhd:3277:73  */
  always @*
    case (n4993)
      2'b10: n5005 = n4978;
      2'b01: n5005 = frestore_fp_temp;
      default: n5005 = frestore_fp_temp;
    endcase
  /* TG68K_FPU.vhd:3275:65  */
  assign n5008 = $unsigned(fsave_counter) >= $unsigned(6'b011100);
  /* TG68K_FPU.vhd:3275:65  */
  assign n5009 = $unsigned(fsave_counter) <= $unsigned(6'b110101);
  /* TG68K_FPU.vhd:3275:65  */
  assign n5010 = n5008 & n5009;
  assign n5011 = {n5010, n4858, n4849, n4820, n4780, n4673, n4667};
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5013 = n4994;
      7'b0100000: n5013 = fpu_done_i;
      7'b0010000: n5013 = n4834;
      7'b0001000: n5013 = n4814;
      7'b0000100: n5013 = fpu_done_i;
      7'b0000010: n5013 = fpu_done_i;
      7'b0000001: n5013 = n4632;
      default: n5013 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5014 = fpu_exception_i;
      7'b0100000: n5014 = fpu_exception_i;
      7'b0010000: n5014 = fpu_exception_i;
      7'b0001000: n5014 = fpu_exception_i;
      7'b0000100: n5014 = fpu_exception_i;
      7'b0000010: n5014 = fpu_exception_i;
      7'b0000001: n5014 = n4634;
      default: n5014 = fpu_exception_i;
    endcase
  assign n5015 = n755[79:0]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5016 = n5015;
      7'b0100000: n5016 = n5015;
      7'b0010000: n5016 = n5015;
      7'b0001000: n5016 = n5015;
      7'b0000100: n5016 = n5015;
      7'b0000010: n5016 = n5015;
      7'b0000001: n5016 = n4636;
      default: n5016 = n5015;
    endcase
  assign n5017 = n755[159:80]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5018 = n5017;
      7'b0100000: n5018 = n5017;
      7'b0010000: n5018 = n5017;
      7'b0001000: n5018 = n5017;
      7'b0000100: n5018 = n5017;
      7'b0000010: n5018 = n5017;
      7'b0000001: n5018 = n4638;
      default: n5018 = n5017;
    endcase
  assign n5019 = n755[239:160]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5020 = n5019;
      7'b0100000: n5020 = n5019;
      7'b0010000: n5020 = n5019;
      7'b0001000: n5020 = n5019;
      7'b0000100: n5020 = n5019;
      7'b0000010: n5020 = n5019;
      7'b0000001: n5020 = n4640;
      default: n5020 = n5019;
    endcase
  assign n5021 = n755[319:240]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5022 = n5021;
      7'b0100000: n5022 = n5021;
      7'b0010000: n5022 = n5021;
      7'b0001000: n5022 = n5021;
      7'b0000100: n5022 = n5021;
      7'b0000010: n5022 = n5021;
      7'b0000001: n5022 = n4642;
      default: n5022 = n5021;
    endcase
  assign n5023 = n755[399:320]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5024 = n5023;
      7'b0100000: n5024 = n5023;
      7'b0010000: n5024 = n5023;
      7'b0001000: n5024 = n5023;
      7'b0000100: n5024 = n5023;
      7'b0000010: n5024 = n5023;
      7'b0000001: n5024 = n4644;
      default: n5024 = n5023;
    endcase
  assign n5025 = n755[479:400]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5026 = n5025;
      7'b0100000: n5026 = n5025;
      7'b0010000: n5026 = n5025;
      7'b0001000: n5026 = n5025;
      7'b0000100: n5026 = n5025;
      7'b0000010: n5026 = n5025;
      7'b0000001: n5026 = n4646;
      default: n5026 = n5025;
    endcase
  assign n5027 = n755[559:480]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5028 = n5027;
      7'b0100000: n5028 = n5027;
      7'b0010000: n5028 = n5027;
      7'b0001000: n5028 = n5027;
      7'b0000100: n5028 = n5027;
      7'b0000010: n5028 = n5027;
      7'b0000001: n5028 = n4648;
      default: n5028 = n5027;
    endcase
  assign n5029 = n755[639:560]; // extract
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5030 = n5029;
      7'b0100000: n5030 = n5029;
      7'b0010000: n5030 = n5029;
      7'b0001000: n5030 = n5029;
      7'b0000100: n5030 = n5029;
      7'b0000010: n5030 = n5029;
      7'b0000001: n5030 = n4650;
      default: n5030 = n5029;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5034 = n4998;
      7'b0100000: n5034 = 1'b0;
      7'b0010000: n5034 = 1'b0;
      7'b0001000: n5034 = 1'b0;
      7'b0000100: n5034 = 1'b0;
      7'b0000010: n5034 = 1'b0;
      7'b0000001: n5034 = 1'b0;
      default: n5034 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5035 = n4999;
      7'b0100000: n5035 = fp_reg_write_addr;
      7'b0010000: n5035 = fp_reg_write_addr;
      7'b0001000: n5035 = fp_reg_write_addr;
      7'b0000100: n5035 = fp_reg_write_addr;
      7'b0000010: n5035 = fp_reg_write_addr;
      7'b0000001: n5035 = fp_reg_write_addr;
      default: n5035 = fp_reg_write_addr;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5036 = n5000;
      7'b0100000: n5036 = fp_reg_write_data;
      7'b0010000: n5036 = fp_reg_write_data;
      7'b0001000: n5036 = fp_reg_write_data;
      7'b0000100: n5036 = fp_reg_write_data;
      7'b0000010: n5036 = fp_reg_write_data;
      7'b0000001: n5036 = fp_reg_write_data;
      default: n5036 = fp_reg_write_data;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5038 = n5002;
      7'b0100000: n5038 = 1'b0;
      7'b0010000: n5038 = 1'b0;
      7'b0001000: n5038 = 1'b0;
      7'b0000100: n5038 = 1'b0;
      7'b0000010: n5038 = 1'b0;
      7'b0000001: n5038 = 1'b0;
      default: n5038 = 1'b0;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5039 = fpcr;
      7'b0100000: n5039 = fpcr;
      7'b0010000: n5039 = fpcr;
      7'b0001000: n5039 = fpcr;
      7'b0000100: n5039 = n4767;
      7'b0000010: n5039 = fpcr;
      7'b0000001: n5039 = n4652;
      default: n5039 = fpcr;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5041 = fpsr;
      7'b0100000: n5041 = fpsr;
      7'b0010000: n5041 = fpsr;
      7'b0001000: n5041 = frestore_data_in;
      7'b0000100: n5041 = fpsr;
      7'b0000010: n5041 = fpsr;
      7'b0000001: n5041 = n4654;
      default: n5041 = fpsr;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5044 = fpiar;
      7'b0100000: n5044 = fpiar;
      7'b0010000: n5044 = fpiar;
      7'b0001000: n5044 = fpiar;
      7'b0000100: n5044 = fpiar;
      7'b0000010: n5044 = frestore_data_in;
      7'b0000001: n5044 = n4656;
      default: n5044 = fpiar;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5045 = fpcr_rounding_mode_valid;
      7'b0100000: n5045 = fpcr_rounding_mode_valid;
      7'b0010000: n5045 = fpcr_rounding_mode_valid;
      7'b0001000: n5045 = fpcr_rounding_mode_valid;
      7'b0000100: n5045 = n4772;
      7'b0000010: n5045 = fpcr_rounding_mode_valid;
      7'b0000001: n5045 = fpcr_rounding_mode_valid;
      default: n5045 = fpcr_rounding_mode_valid;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5046 = fpcr_precision_valid;
      7'b0100000: n5046 = fpcr_precision_valid;
      7'b0010000: n5046 = fpcr_precision_valid;
      7'b0001000: n5046 = fpcr_precision_valid;
      7'b0000100: n5046 = n4774;
      7'b0000010: n5046 = fpcr_precision_valid;
      7'b0000001: n5046 = fpcr_precision_valid;
      default: n5046 = fpcr_precision_valid;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5050 = n5003;
      7'b0100000: n5050 = fpu_state;
      7'b0010000: n5050 = n4836;
      7'b0001000: n5050 = n4817;
      7'b0000100: n5050 = fpu_state;
      7'b0000010: n5050 = fpu_state;
      7'b0000001: n5050 = n4660;
      default: n5050 = 4'b0000;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5051 = fpu_just_reset;
      7'b0100000: n5051 = fpu_just_reset;
      7'b0010000: n5051 = fpu_just_reset;
      7'b0001000: n5051 = fpu_just_reset;
      7'b0000100: n5051 = fpu_just_reset;
      7'b0000010: n5051 = fpu_just_reset;
      7'b0000001: n5051 = n4662;
      default: n5051 = fpu_just_reset;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5052 = n5004;
      7'b0100000: n5052 = n4853;
      7'b0010000: n5052 = n4844;
      7'b0001000: n5052 = n4818;
      7'b0000100: n5052 = n4778;
      7'b0000010: n5052 = n4671;
      7'b0000001: n5052 = n4663;
      default: n5052 = fsave_counter;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5053 = frestore_frame_format;
      7'b0100000: n5053 = frestore_frame_format;
      7'b0010000: n5053 = frestore_frame_format;
      7'b0001000: n5053 = frestore_frame_format;
      7'b0000100: n5053 = frestore_frame_format;
      7'b0000010: n5053 = frestore_frame_format;
      7'b0000001: n5053 = n4591;
      default: n5053 = frestore_frame_format;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5054 = n5005;
      7'b0100000: n5054 = frestore_fp_temp;
      7'b0010000: n5054 = frestore_fp_temp;
      7'b0001000: n5054 = frestore_fp_temp;
      7'b0000100: n5054 = frestore_fp_temp;
      7'b0000010: n5054 = frestore_fp_temp;
      7'b0000001: n5054 = frestore_fp_temp;
      default: n5054 = frestore_fp_temp;
    endcase
  /* TG68K_FPU.vhd:3147:57  */
  always @*
    case (n5011)
      7'b1000000: n5055 = exception_code_internal;
      7'b0100000: n5055 = exception_code_internal;
      7'b0010000: n5055 = exception_code_internal;
      7'b0001000: n5055 = exception_code_internal;
      7'b0000100: n5055 = exception_code_internal;
      7'b0000010: n5055 = exception_code_internal;
      7'b0000001: n5055 = n4665;
      default: n5055 = exception_code_internal;
    endcase
  /* TG68K_FPU.vhd:3145:49  */
  assign n5056 = frestore_data_write ? n5013 : fpu_done_i;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5057 = frestore_data_write ? n5014 : fpu_exception_i;
  assign n5058 = {n5030, n5028, n5026, n5024, n5022, n5020, n5018, n5016};
  /* TG68K_FPU.vhd:3145:49  */
  assign n5059 = frestore_data_write ? n5058 : n755;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5063 = frestore_data_write ? n5034 : 1'b0;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5065 = frestore_data_write ? n5035 : fp_reg_write_addr;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5066 = frestore_data_write ? n5036 : fp_reg_write_data;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5068 = frestore_data_write ? n5038 : 1'b0;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5070 = frestore_data_write ? n5039 : fpcr;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5072 = frestore_data_write ? n5041 : fpsr;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5074 = frestore_data_write ? n5044 : fpiar;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5075 = frestore_data_write ? n5045 : fpcr_rounding_mode_valid;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5076 = frestore_data_write ? n5046 : fpcr_precision_valid;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5078 = frestore_data_write ? n5050 : fpu_state;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5079 = frestore_data_write ? n5051 : fpu_just_reset;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5080 = frestore_data_write ? n5052 : fsave_counter;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5081 = frestore_data_write ? n5053 : frestore_frame_format;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5082 = frestore_data_write ? n5054 : frestore_fp_temp;
  /* TG68K_FPU.vhd:3145:49  */
  assign n5083 = frestore_data_write ? n5055 : exception_code_internal;
  /* TG68K_FPU.vhd:3139:41  */
  assign n5085 = fpu_state == 4'b1010;
  /* TG68K_FPU.vhd:3358:65  */
  assign n5088 = fmovem_reg_index == 3'b000;
  /* TG68K_FPU.vhd:3367:65  */
  assign n5091 = fmovem_reg_index == 3'b001;
  /* TG68K_FPU.vhd:3376:65  */
  assign n5094 = fmovem_reg_index == 3'b010;
  /* TG68K_FPU.vhd:3385:65  */
  assign n5097 = fmovem_reg_index == 3'b011;
  /* TG68K_FPU.vhd:3394:65  */
  assign n5100 = fmovem_reg_index == 3'b100;
  /* TG68K_FPU.vhd:3403:65  */
  assign n5103 = fmovem_reg_index == 3'b101;
  /* TG68K_FPU.vhd:3412:65  */
  assign n5106 = fmovem_reg_index == 3'b110;
  /* TG68K_FPU.vhd:3421:65  */
  assign n5109 = fmovem_reg_index == 3'b111;
  assign n5110 = {n5109, n5106, n5103, n5100, n5097, n5094, n5091, n5088};
  /* TG68K_FPU.vhd:3357:57  */
  always @*
    case (n5110)
      8'b10000000: n5144 = 1'b1;
      8'b01000000: n5144 = 1'b1;
      8'b00100000: n5144 = 1'b1;
      8'b00010000: n5144 = 1'b1;
      8'b00001000: n5144 = 1'b1;
      8'b00000100: n5144 = 1'b1;
      8'b00000010: n5144 = 1'b1;
      8'b00000001: n5144 = 1'b1;
      default: n5144 = fp_reg_write_enable;
    endcase
  /* TG68K_FPU.vhd:3357:57  */
  always @*
    case (n5110)
      8'b10000000: n5153 = 3'b111;
      8'b01000000: n5153 = 3'b110;
      8'b00100000: n5153 = 3'b101;
      8'b00010000: n5153 = 3'b100;
      8'b00001000: n5153 = 3'b011;
      8'b00000100: n5153 = 3'b010;
      8'b00000010: n5153 = 3'b001;
      8'b00000001: n5153 = 3'b000;
      default: n5153 = fp_reg_write_addr;
    endcase
  /* TG68K_FPU.vhd:3357:57  */
  always @*
    case (n5110)
      8'b10000000: n5154 = fmovem_data_in;
      8'b01000000: n5154 = fmovem_data_in;
      8'b00100000: n5154 = fmovem_data_in;
      8'b00010000: n5154 = fmovem_data_in;
      8'b00001000: n5154 = fmovem_data_in;
      8'b00000100: n5154 = fmovem_data_in;
      8'b00000010: n5154 = fmovem_data_in;
      8'b00000001: n5154 = fmovem_data_in;
      default: n5154 = fp_reg_write_data;
    endcase
  /* TG68K_FPU.vhd:3357:57  */
  always @*
    case (n5110)
      8'b10000000: n5163 = 1'b1;
      8'b01000000: n5163 = 1'b1;
      8'b00100000: n5163 = 1'b1;
      8'b00010000: n5163 = 1'b1;
      8'b00001000: n5163 = 1'b1;
      8'b00000100: n5163 = 1'b1;
      8'b00000010: n5163 = 1'b1;
      8'b00000001: n5163 = 1'b1;
      default: n5163 = fp_reg_access_valid;
    endcase
  /* TG68K_FPU.vhd:3354:49  */
  assign n5167 = fmovem_data_write ? n5144 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:3354:49  */
  assign n5168 = fmovem_data_write ? n5153 : fp_reg_write_addr;
  /* TG68K_FPU.vhd:3354:49  */
  assign n5169 = fmovem_data_write ? n5154 : fp_reg_write_data;
  /* TG68K_FPU.vhd:3354:49  */
  assign n5170 = fmovem_data_write ? n5163 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:3437:63  */
  assign n5171 = ~fpu_enable;
  /* TG68K_FPU.vhd:3437:69  */
  assign n5172 = n5171 | movem_done;
  /* TG68K_FPU.vhd:3437:49  */
  assign n5174 = n5172 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3437:49  */
  assign n5176 = n5172 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3346:41  */
  assign n5178 = fpu_state == 4'b1011;
  /* TG68K_FPU.vhd:3449:65  */
  assign n5180 = fmovem_reg_index == 3'b000;
  /* TG68K_FPU.vhd:3450:65  */
  assign n5182 = fmovem_reg_index == 3'b001;
  /* TG68K_FPU.vhd:3451:65  */
  assign n5184 = fmovem_reg_index == 3'b010;
  assign n5185 = {n5184, n5182, n5180};
  /* TG68K_FPU.vhd:3448:57  */
  always @*
    case (n5185)
      3'b100: n5187 = fpiar;
      3'b010: n5187 = fpsr;
      3'b001: n5187 = fpcr;
      default: n5187 = 32'b00000000000000000000000000000000;
    endcase
  /* TG68K_FPU.vhd:3447:49  */
  assign n5188 = fmovem_data_request ? n5187 : n6841;
  /* TG68K_FPU.vhd:613:28  */
  assign n5194 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:613:41  */
  assign n5196 = n5194 == 2'b11;
  /* TG68K_FPU.vhd:613:17  */
  assign n5200 = n5196 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:613:17  */
  assign n5206 = n5196 ? 1'b0 : 1'bX;
  /* TG68K_FPU.vhd:618:28  */
  assign n5207 = cpu_data_in[31:16]; // extract
  /* TG68K_FPU.vhd:618:43  */
  assign n5209 = n5207 != 16'b0000000000000000;
  /* TG68K_FPU.vhd:618:65  */
  assign n5210 = cpu_data_in[5:0]; // extract
  /* TG68K_FPU.vhd:618:78  */
  assign n5212 = n5210 != 6'b000000;
  /* TG68K_FPU.vhd:618:54  */
  assign n5213 = n5209 | n5212;
  /* TG68K_FPU.vhd:618:17  */
  assign n5216 = n5223 ? 1'b0 : n5200;
  /* TG68K_FPU.vhd:618:17  */
  assign n5219 = n5225 ? 1'b0 : n5206;
  /* TG68K_FPU.vhd:618:17  */
  assign n5220 = n5200 & n5213;
  /* TG68K_FPU.vhd:618:17  */
  assign n5222 = n5200 & n5213;
  /* TG68K_FPU.vhd:618:17  */
  assign n5223 = n5220 & n5200;
  /* TG68K_FPU.vhd:618:17  */
  assign n5225 = n5222 & n5200;
  /* TG68K_FPU.vhd:623:17  */
  assign n5231 = n5216 ? 1'b1 : n5219;
  /* TG68K_FPU.vhd:597:30  */
  assign n5239 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:43  */
  assign n5241 = n5239 == 2'b11;
  assign n5243 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:17  */
  assign n5244 = n5241 ? 2'b00 : n5243;
  assign n5248 = cpu_data_in[15:8]; // extract
  assign n5250 = {16'b0000000000000000, n5248, n5244, 6'b000000};
  /* TG68K_FPU.vhd:597:30  */
  assign n5258 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:43  */
  assign n5260 = n5258 == 2'b11;
  assign n5262 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:597:17  */
  assign n5263 = n5260 ? 2'b00 : n5262;
  assign n5267 = cpu_data_in[15:8]; // extract
  assign n5269 = {16'b0000000000000000, n5267, n5263, 6'b000000};
  /* TG68K_FPU.vhd:3470:95  */
  assign n5270 = cpu_data_in[15:14]; // extract
  /* TG68K_FPU.vhd:3470:110  */
  assign n5272 = n5270 == 2'b11;
  /* TG68K_FPU.vhd:3470:81  */
  assign n5275 = n5272 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:3475:95  */
  assign n5276 = cpu_data_in[7:6]; // extract
  /* TG68K_FPU.vhd:3475:108  */
  assign n5278 = n5276 == 2'b11;
  /* TG68K_FPU.vhd:3475:81  */
  assign n5281 = n5278 ? 1'b0 : 1'b1;
  /* TG68K_FPU.vhd:3461:73  */
  assign n5282 = n5231 ? n5250 : n5269;
  /* TG68K_FPU.vhd:3461:73  */
  assign n5287 = n5231 ? 1'b1 : n5275;
  /* TG68K_FPU.vhd:3461:73  */
  assign n5289 = n5231 ? 1'b1 : n5281;
  /* TG68K_FPU.vhd:3459:65  */
  assign n5291 = fmovem_reg_index == 3'b000;
  /* TG68K_FPU.vhd:3481:65  */
  assign n5300 = fmovem_reg_index == 3'b001;
  /* TG68K_FPU.vhd:3486:65  */
  assign n5302 = fmovem_reg_index == 3'b010;
  assign n5303 = {n5302, n5300, n5291};
  /* TG68K_FPU.vhd:3458:57  */
  always @*
    case (n5303)
      3'b100: n5304 = fpcr;
      3'b010: n5304 = fpcr;
      3'b001: n5304 = n5282;
      default: n5304 = fpcr;
    endcase
  /* TG68K_FPU.vhd:3458:57  */
  always @*
    case (n5303)
      3'b100: n5306 = fpsr;
      3'b010: n5306 = cpu_data_in;
      3'b001: n5306 = fpsr;
      default: n5306 = fpsr;
    endcase
  /* TG68K_FPU.vhd:3458:57  */
  always @*
    case (n5303)
      3'b100: n5309 = cpu_data_in;
      3'b010: n5309 = fpiar;
      3'b001: n5309 = fpiar;
      default: n5309 = fpiar;
    endcase
  /* TG68K_FPU.vhd:3458:57  */
  always @*
    case (n5303)
      3'b100: n5312 = fpcr_rounding_mode_valid;
      3'b010: n5312 = fpcr_rounding_mode_valid;
      3'b001: n5312 = n5287;
      default: n5312 = fpcr_rounding_mode_valid;
    endcase
  /* TG68K_FPU.vhd:3458:57  */
  always @*
    case (n5303)
      3'b100: n5313 = fpcr_precision_valid;
      3'b010: n5313 = fpcr_precision_valid;
      3'b001: n5313 = n5289;
      default: n5313 = fpcr_precision_valid;
    endcase
  /* TG68K_FPU.vhd:3457:49  */
  assign n5316 = fmovem_data_write ? n5304 : fpcr;
  /* TG68K_FPU.vhd:3457:49  */
  assign n5318 = fmovem_data_write ? n5306 : fpsr;
  /* TG68K_FPU.vhd:3457:49  */
  assign n5320 = fmovem_data_write ? n5309 : fpiar;
  /* TG68K_FPU.vhd:3457:49  */
  assign n5322 = fmovem_data_write ? n5312 : fpcr_rounding_mode_valid;
  /* TG68K_FPU.vhd:3457:49  */
  assign n5323 = fmovem_data_write ? n5313 : fpcr_precision_valid;
  /* TG68K_FPU.vhd:3495:63  */
  assign n5325 = ~fpu_enable;
  /* TG68K_FPU.vhd:3495:69  */
  assign n5326 = n5325 | movem_done;
  /* TG68K_FPU.vhd:3495:49  */
  assign n5328 = n5326 ? 1'b1 : fpu_done_i;
  /* TG68K_FPU.vhd:3495:49  */
  assign n5330 = n5326 ? 4'b0000 : fpu_state;
  /* TG68K_FPU.vhd:3442:41  */
  assign n5332 = fpu_state == 4'b1100;
  assign n5333 = {n5332, n5178, n5085, n4590, n4448, n4350, n4348, n4047, n4045, n4043, n3643, n2790, n855};
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5337 = n5188;
      13'b0100000000000: n5337 = n6841;
      13'b0010000000000: n5337 = n6841;
      13'b0001000000000: n5337 = n4547;
      13'b0000100000000: n5337 = n6841;
      13'b0000010000000: n5337 = n6841;
      13'b0000001000000: n5337 = n4327;
      13'b0000000100000: n5337 = n6841;
      13'b0000000010000: n5337 = n6841;
      13'b0000000001000: n5337 = 32'b00000000000000000000000000000000;
      13'b0000000000100: n5337 = 32'b00000000000000000000000000000000;
      13'b0000000000010: n5337 = n2750;
      13'b0000000000001: n5337 = n841;
      default: n5337 = 32'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5342 = n5328;
      13'b0100000000000: n5342 = n5174;
      13'b0010000000000: n5342 = n5056;
      13'b0001000000000: n5342 = n4587;
      13'b0000100000000: n5342 = 1'b1;
      13'b0000010000000: n5342 = 1'b1;
      13'b0000001000000: n5342 = n4329;
      13'b0000000100000: n5342 = 1'b1;
      13'b0000000010000: n5342 = fpu_done_i;
      13'b0000000001000: n5342 = n4026;
      13'b0000000000100: n5342 = fpu_done_i;
      13'b0000000000010: n5342 = n2753;
      13'b0000000000001: n5342 = n843;
      default: n5342 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5344 = fpu_exception_i;
      13'b0100000000000: n5344 = fpu_exception_i;
      13'b0010000000000: n5344 = n5057;
      13'b0001000000000: n5344 = fpu_exception_i;
      13'b0000100000000: n5344 = n4446;
      13'b0000010000000: n5344 = fpu_exception_i;
      13'b0000001000000: n5344 = n4068;
      13'b0000000100000: n5344 = fpu_exception_i;
      13'b0000000010000: n5344 = fpu_exception_i;
      13'b0000000001000: n5344 = n4027;
      13'b0000000000100: n5344 = n3626;
      13'b0000000000010: n5344 = n2755;
      13'b0000000000001: n5344 = n844;
      default: n5344 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5346 = n755;
      13'b0100000000000: n5346 = n755;
      13'b0010000000000: n5346 = n5059;
      13'b0001000000000: n5346 = n755;
      13'b0000100000000: n5346 = n755;
      13'b0000010000000: n5346 = n755;
      13'b0000001000000: n5346 = n755;
      13'b0000000100000: n5346 = n755;
      13'b0000000010000: n5346 = n755;
      13'b0000000001000: n5346 = n755;
      13'b0000000000100: n5346 = n755;
      13'b0000000000010: n5346 = n755;
      13'b0000000000001: n5346 = n755;
      default: n5346 = 640'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5352 = fp_reg_write_enable;
      13'b0100000000000: n5352 = n5167;
      13'b0010000000000: n5352 = n5063;
      13'b0001000000000: n5352 = fp_reg_write_enable;
      13'b0000100000000: n5352 = fp_reg_write_enable;
      13'b0000010000000: n5352 = fp_reg_write_enable;
      13'b0000001000000: n5352 = n4333;
      13'b0000000100000: n5352 = fp_reg_write_enable;
      13'b0000000010000: n5352 = fp_reg_write_enable;
      13'b0000000001000: n5352 = fp_reg_write_enable;
      13'b0000000000100: n5352 = fp_reg_write_enable;
      13'b0000000000010: n5352 = n2756;
      13'b0000000000001: n5352 = fp_reg_write_enable;
      default: n5352 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5354 = fp_reg_write_addr;
      13'b0100000000000: n5354 = n5168;
      13'b0010000000000: n5354 = n5065;
      13'b0001000000000: n5354 = fp_reg_write_addr;
      13'b0000100000000: n5354 = fp_reg_write_addr;
      13'b0000010000000: n5354 = fp_reg_write_addr;
      13'b0000001000000: n5354 = n4334;
      13'b0000000100000: n5354 = fp_reg_write_addr;
      13'b0000000010000: n5354 = fp_reg_write_addr;
      13'b0000000001000: n5354 = fp_reg_write_addr;
      13'b0000000000100: n5354 = fp_reg_write_addr;
      13'b0000000000010: n5354 = n2757;
      13'b0000000000001: n5354 = fp_reg_write_addr;
      default: n5354 = 3'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5356 = fp_reg_write_data;
      13'b0100000000000: n5356 = n5169;
      13'b0010000000000: n5356 = n5066;
      13'b0001000000000: n5356 = fp_reg_write_data;
      13'b0000100000000: n5356 = fp_reg_write_data;
      13'b0000010000000: n5356 = fp_reg_write_data;
      13'b0000001000000: n5356 = n4335;
      13'b0000000100000: n5356 = fp_reg_write_data;
      13'b0000000010000: n5356 = fp_reg_write_data;
      13'b0000000001000: n5356 = fp_reg_write_data;
      13'b0000000000100: n5356 = fp_reg_write_data;
      13'b0000000000010: n5356 = n2758;
      13'b0000000000001: n5356 = fp_reg_write_data;
      default: n5356 = 80'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5360 = fp_reg_access_valid;
      13'b0100000000000: n5360 = n5170;
      13'b0010000000000: n5360 = n5068;
      13'b0001000000000: n5360 = fp_reg_access_valid;
      13'b0000100000000: n5360 = fp_reg_access_valid;
      13'b0000010000000: n5360 = fp_reg_access_valid;
      13'b0000001000000: n5360 = n4336;
      13'b0000000100000: n5360 = fp_reg_access_valid;
      13'b0000000010000: n5360 = fp_reg_access_valid;
      13'b0000000001000: n5360 = fp_reg_access_valid;
      13'b0000000000100: n5360 = fp_reg_access_valid;
      13'b0000000000010: n5360 = n2760;
      13'b0000000000001: n5360 = fp_reg_access_valid;
      default: n5360 = 1'bX;
    endcase
  assign n5361 = n2761[5:0]; // extract
  assign n5362 = n5070[5:0]; // extract
  assign n5363 = n5316[5:0]; // extract
  assign n5364 = fpcr[5:0]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5366 = n5363;
      13'b0100000000000: n5366 = n5364;
      13'b0010000000000: n5366 = n5362;
      13'b0001000000000: n5366 = n5364;
      13'b0000100000000: n5366 = n5364;
      13'b0000010000000: n5366 = n5364;
      13'b0000001000000: n5366 = n5364;
      13'b0000000100000: n5366 = n5364;
      13'b0000000010000: n5366 = n5364;
      13'b0000000001000: n5366 = n5364;
      13'b0000000000100: n5366 = n5364;
      13'b0000000000010: n5366 = n5361;
      13'b0000000000001: n5366 = n5364;
      default: n5366 = 6'bX;
    endcase
  assign n5367 = n2761[7:6]; // extract
  assign n5368 = n5070[7:6]; // extract
  assign n5369 = n5316[7:6]; // extract
  assign n5370 = fpcr[7:6]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5372 = n5369;
      13'b0100000000000: n5372 = n5370;
      13'b0010000000000: n5372 = n5368;
      13'b0001000000000: n5372 = n5370;
      13'b0000100000000: n5372 = n5370;
      13'b0000010000000: n5372 = n5370;
      13'b0000001000000: n5372 = n5370;
      13'b0000000100000: n5372 = n5370;
      13'b0000000010000: n5372 = n5370;
      13'b0000000001000: n5372 = n3681;
      13'b0000000000100: n5372 = n5370;
      13'b0000000000010: n5372 = n5367;
      13'b0000000000001: n5372 = n5370;
      default: n5372 = 2'bX;
    endcase
  assign n5373 = n2761[13:8]; // extract
  assign n5374 = n5070[13:8]; // extract
  assign n5375 = n5316[13:8]; // extract
  assign n5376 = fpcr[13:8]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5378 = n5375;
      13'b0100000000000: n5378 = n5376;
      13'b0010000000000: n5378 = n5374;
      13'b0001000000000: n5378 = n5376;
      13'b0000100000000: n5378 = n5376;
      13'b0000010000000: n5378 = n5376;
      13'b0000001000000: n5378 = n5376;
      13'b0000000100000: n5378 = n5376;
      13'b0000000010000: n5378 = n5376;
      13'b0000000001000: n5378 = n5376;
      13'b0000000000100: n5378 = n5376;
      13'b0000000000010: n5378 = n5373;
      13'b0000000000001: n5378 = n5376;
      default: n5378 = 6'bX;
    endcase
  assign n5379 = n2761[15:14]; // extract
  assign n5380 = n5070[15:14]; // extract
  assign n5381 = n5316[15:14]; // extract
  assign n5382 = fpcr[15:14]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5384 = n5381;
      13'b0100000000000: n5384 = n5382;
      13'b0010000000000: n5384 = n5380;
      13'b0001000000000: n5384 = n5382;
      13'b0000100000000: n5384 = n5382;
      13'b0000010000000: n5384 = n5382;
      13'b0000001000000: n5384 = n5382;
      13'b0000000100000: n5384 = n5382;
      13'b0000000010000: n5384 = n5382;
      13'b0000000001000: n5384 = n3663;
      13'b0000000000100: n5384 = n5382;
      13'b0000000000010: n5384 = n5379;
      13'b0000000000001: n5384 = n5382;
      default: n5384 = 2'bX;
    endcase
  assign n5385 = n2761[31:16]; // extract
  assign n5386 = n5070[31:16]; // extract
  assign n5387 = n5316[31:16]; // extract
  assign n5388 = fpcr[31:16]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5390 = n5387;
      13'b0100000000000: n5390 = n5388;
      13'b0010000000000: n5390 = n5386;
      13'b0001000000000: n5390 = n5388;
      13'b0000100000000: n5390 = n5388;
      13'b0000010000000: n5390 = n5388;
      13'b0000001000000: n5390 = n5388;
      13'b0000000100000: n5390 = n5388;
      13'b0000000010000: n5390 = n5388;
      13'b0000000001000: n5390 = n5388;
      13'b0000000000100: n5390 = n5388;
      13'b0000000000010: n5390 = n5385;
      13'b0000000000001: n5390 = n5388;
      default: n5390 = 16'bX;
    endcase
  assign n5395 = n2762[12:0]; // extract
  assign n5396 = n4028[12:0]; // extract
  assign n5397 = n5072[12:0]; // extract
  assign n5398 = n5318[12:0]; // extract
  assign n5399 = fpsr[12:0]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5401 = n5398;
      13'b0100000000000: n5401 = n5399;
      13'b0010000000000: n5401 = n5397;
      13'b0001000000000: n5401 = n5399;
      13'b0000100000000: n5401 = n5399;
      13'b0000010000000: n5401 = n5399;
      13'b0000001000000: n5401 = n5399;
      13'b0000000100000: n5401 = n5399;
      13'b0000000010000: n5401 = n5399;
      13'b0000000001000: n5401 = n5396;
      13'b0000000000100: n5401 = n5399;
      13'b0000000000010: n5401 = n5395;
      13'b0000000000001: n5401 = n5399;
      default: n5401 = 13'bX;
    endcase
  assign n5402 = n2762[13]; // extract
  assign n5403 = n4028[13]; // extract
  assign n5404 = n5072[13]; // extract
  assign n5405 = n5318[13]; // extract
  assign n5406 = fpsr[13]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5408 = n5405;
      13'b0100000000000: n5408 = n5406;
      13'b0010000000000: n5408 = n5404;
      13'b0001000000000: n5408 = n5406;
      13'b0000100000000: n5408 = n4385;
      13'b0000010000000: n5408 = n5406;
      13'b0000001000000: n5408 = n5406;
      13'b0000000100000: n5408 = n5406;
      13'b0000000010000: n5408 = n5406;
      13'b0000000001000: n5408 = n5403;
      13'b0000000000100: n5408 = n5406;
      13'b0000000000010: n5408 = n5402;
      13'b0000000000001: n5408 = n5406;
      default: n5408 = 1'bX;
    endcase
  assign n5409 = n2762[14]; // extract
  assign n5410 = n4028[14]; // extract
  assign n5411 = n4340[0]; // extract
  assign n5412 = n5072[14]; // extract
  assign n5413 = n5318[14]; // extract
  assign n5414 = fpsr[14]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5416 = n5413;
      13'b0100000000000: n5416 = n5414;
      13'b0010000000000: n5416 = n5412;
      13'b0001000000000: n5416 = n5414;
      13'b0000100000000: n5416 = n4387;
      13'b0000010000000: n5416 = n5414;
      13'b0000001000000: n5416 = n5411;
      13'b0000000100000: n5416 = n5414;
      13'b0000000010000: n5416 = n5414;
      13'b0000000001000: n5416 = n5410;
      13'b0000000000100: n5416 = n5414;
      13'b0000000000010: n5416 = n5409;
      13'b0000000000001: n5416 = n5414;
      default: n5416 = 1'bX;
    endcase
  assign n5417 = n2762[15]; // extract
  assign n5418 = n4028[15]; // extract
  assign n5419 = n4340[1]; // extract
  assign n5420 = n5072[15]; // extract
  assign n5421 = n5318[15]; // extract
  assign n5422 = fpsr[15]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5424 = n5421;
      13'b0100000000000: n5424 = n5422;
      13'b0010000000000: n5424 = n5420;
      13'b0001000000000: n5424 = n5422;
      13'b0000100000000: n5424 = n4389;
      13'b0000010000000: n5424 = n5422;
      13'b0000001000000: n5424 = n5419;
      13'b0000000100000: n5424 = n5422;
      13'b0000000010000: n5424 = n5422;
      13'b0000000001000: n5424 = n5418;
      13'b0000000000100: n5424 = n5422;
      13'b0000000000010: n5424 = n5417;
      13'b0000000000001: n5424 = n5422;
      default: n5424 = 1'bX;
    endcase
  assign n5425 = n2762[16]; // extract
  assign n5426 = n4028[16]; // extract
  assign n5427 = n4340[2]; // extract
  assign n5428 = n5072[16]; // extract
  assign n5429 = n5318[16]; // extract
  assign n5430 = fpsr[16]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5432 = n5429;
      13'b0100000000000: n5432 = n5430;
      13'b0010000000000: n5432 = n5428;
      13'b0001000000000: n5432 = n5430;
      13'b0000100000000: n5432 = n4391;
      13'b0000010000000: n5432 = n5430;
      13'b0000001000000: n5432 = n5427;
      13'b0000000100000: n5432 = n5430;
      13'b0000000010000: n5432 = n5430;
      13'b0000000001000: n5432 = n5426;
      13'b0000000000100: n5432 = n5430;
      13'b0000000000010: n5432 = n5425;
      13'b0000000000001: n5432 = n5430;
      default: n5432 = 1'bX;
    endcase
  assign n5433 = n2762[17]; // extract
  assign n5434 = n4028[17]; // extract
  assign n5435 = n4340[3]; // extract
  assign n5436 = n5072[17]; // extract
  assign n5437 = n5318[17]; // extract
  assign n5438 = fpsr[17]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5440 = n5437;
      13'b0100000000000: n5440 = n5438;
      13'b0010000000000: n5440 = n5436;
      13'b0001000000000: n5440 = n5438;
      13'b0000100000000: n5440 = n4393;
      13'b0000010000000: n5440 = n5438;
      13'b0000001000000: n5440 = n5435;
      13'b0000000100000: n5440 = n5438;
      13'b0000000010000: n5440 = n5438;
      13'b0000000001000: n5440 = n5434;
      13'b0000000000100: n5440 = n5438;
      13'b0000000000010: n5440 = n5433;
      13'b0000000000001: n5440 = n5438;
      default: n5440 = 1'bX;
    endcase
  assign n5441 = n2762[18]; // extract
  assign n5442 = n4028[18]; // extract
  assign n5443 = n4340[4]; // extract
  assign n5444 = n5072[18]; // extract
  assign n5445 = n5318[18]; // extract
  assign n5446 = fpsr[18]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5448 = n5445;
      13'b0100000000000: n5448 = n5446;
      13'b0010000000000: n5448 = n5444;
      13'b0001000000000: n5448 = n5446;
      13'b0000100000000: n5448 = n4395;
      13'b0000010000000: n5448 = n5446;
      13'b0000001000000: n5448 = n5443;
      13'b0000000100000: n5448 = n5446;
      13'b0000000010000: n5448 = n5446;
      13'b0000000001000: n5448 = n5442;
      13'b0000000000100: n5448 = n5446;
      13'b0000000000010: n5448 = n5441;
      13'b0000000000001: n5448 = n5446;
      default: n5448 = 1'bX;
    endcase
  assign n5449 = n2762[20:19]; // extract
  assign n5450 = n4028[20:19]; // extract
  assign n5451 = n4340[6:5]; // extract
  assign n5452 = n5072[20:19]; // extract
  assign n5453 = n5318[20:19]; // extract
  assign n5454 = fpsr[20:19]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5456 = n5453;
      13'b0100000000000: n5456 = n5454;
      13'b0010000000000: n5456 = n5452;
      13'b0001000000000: n5456 = n5454;
      13'b0000100000000: n5456 = n5454;
      13'b0000010000000: n5456 = n5454;
      13'b0000001000000: n5456 = n5451;
      13'b0000000100000: n5456 = n5454;
      13'b0000000010000: n5456 = n5454;
      13'b0000000001000: n5456 = n5450;
      13'b0000000000100: n5456 = n5454;
      13'b0000000000010: n5456 = n5449;
      13'b0000000000001: n5456 = n5454;
      default: n5456 = 2'bX;
    endcase
  assign n5457 = n2762[21]; // extract
  assign n5458 = n4028[21]; // extract
  assign n5459 = n4340[7]; // extract
  assign n5460 = n5072[21]; // extract
  assign n5461 = n5318[21]; // extract
  assign n5462 = fpsr[21]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5464 = n5461;
      13'b0100000000000: n5464 = n5462;
      13'b0010000000000: n5464 = n5460;
      13'b0001000000000: n5464 = n5462;
      13'b0000100000000: n5464 = n4397;
      13'b0000010000000: n5464 = n5462;
      13'b0000001000000: n5464 = n5459;
      13'b0000000100000: n5464 = n5462;
      13'b0000000010000: n5464 = n5462;
      13'b0000000001000: n5464 = n5458;
      13'b0000000000100: n5464 = n5462;
      13'b0000000000010: n5464 = n5457;
      13'b0000000000001: n5464 = n5462;
      default: n5464 = 1'bX;
    endcase
  assign n5465 = n2762[22]; // extract
  assign n5466 = n4028[22]; // extract
  assign n5467 = n4340[8]; // extract
  assign n5468 = n5072[22]; // extract
  assign n5469 = n5318[22]; // extract
  assign n5470 = fpsr[22]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5472 = n5469;
      13'b0100000000000: n5472 = n5470;
      13'b0010000000000: n5472 = n5468;
      13'b0001000000000: n5472 = n5470;
      13'b0000100000000: n5472 = n4399;
      13'b0000010000000: n5472 = n5470;
      13'b0000001000000: n5472 = n5467;
      13'b0000000100000: n5472 = n5470;
      13'b0000000010000: n5472 = n5470;
      13'b0000000001000: n5472 = n5466;
      13'b0000000000100: n5472 = n5470;
      13'b0000000000010: n5472 = n5465;
      13'b0000000000001: n5472 = n5470;
      default: n5472 = 1'bX;
    endcase
  assign n5473 = n2762[23]; // extract
  assign n5474 = n4028[23]; // extract
  assign n5475 = n4340[9]; // extract
  assign n5476 = n5072[23]; // extract
  assign n5477 = n5318[23]; // extract
  assign n5478 = fpsr[23]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5480 = n5477;
      13'b0100000000000: n5480 = n5478;
      13'b0010000000000: n5480 = n5476;
      13'b0001000000000: n5480 = n5478;
      13'b0000100000000: n5480 = n4401;
      13'b0000010000000: n5480 = n5478;
      13'b0000001000000: n5480 = n5475;
      13'b0000000100000: n5480 = n5478;
      13'b0000000010000: n5480 = n5478;
      13'b0000000001000: n5480 = n5474;
      13'b0000000000100: n5480 = n5478;
      13'b0000000000010: n5480 = n5473;
      13'b0000000000001: n5480 = n5478;
      default: n5480 = 1'bX;
    endcase
  assign n5481 = n2762[24]; // extract
  assign n5482 = n4028[24]; // extract
  assign n5483 = n4340[10]; // extract
  assign n5484 = n5072[24]; // extract
  assign n5485 = n5318[24]; // extract
  assign n5486 = fpsr[24]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5488 = n5485;
      13'b0100000000000: n5488 = n5486;
      13'b0010000000000: n5488 = n5484;
      13'b0001000000000: n5488 = n5486;
      13'b0000100000000: n5488 = n4403;
      13'b0000010000000: n5488 = n5486;
      13'b0000001000000: n5488 = n5483;
      13'b0000000100000: n5488 = n5486;
      13'b0000000010000: n5488 = n5486;
      13'b0000000001000: n5488 = n5482;
      13'b0000000000100: n5488 = n5486;
      13'b0000000000010: n5488 = n5481;
      13'b0000000000001: n5488 = n5486;
      default: n5488 = 1'bX;
    endcase
  assign n5489 = n2762[25]; // extract
  assign n5490 = n4028[25]; // extract
  assign n5491 = n4340[11]; // extract
  assign n5492 = n5072[25]; // extract
  assign n5493 = n5318[25]; // extract
  assign n5494 = fpsr[25]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5496 = n5493;
      13'b0100000000000: n5496 = n5494;
      13'b0010000000000: n5496 = n5492;
      13'b0001000000000: n5496 = n5494;
      13'b0000100000000: n5496 = n4405;
      13'b0000010000000: n5496 = n5494;
      13'b0000001000000: n5496 = n5491;
      13'b0000000100000: n5496 = n5494;
      13'b0000000010000: n5496 = n5494;
      13'b0000000001000: n5496 = n5490;
      13'b0000000000100: n5496 = n5494;
      13'b0000000000010: n5496 = n5489;
      13'b0000000000001: n5496 = n5494;
      default: n5496 = 1'bX;
    endcase
  assign n5497 = n2762[26]; // extract
  assign n5498 = n4028[26]; // extract
  assign n5499 = n4340[12]; // extract
  assign n5500 = n5072[26]; // extract
  assign n5501 = n5318[26]; // extract
  assign n5502 = fpsr[26]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5504 = n5501;
      13'b0100000000000: n5504 = n5502;
      13'b0010000000000: n5504 = n5500;
      13'b0001000000000: n5504 = n5502;
      13'b0000100000000: n5504 = n4407;
      13'b0000010000000: n5504 = n5502;
      13'b0000001000000: n5504 = n5499;
      13'b0000000100000: n5504 = n5502;
      13'b0000000010000: n5504 = n5502;
      13'b0000000001000: n5504 = n5498;
      13'b0000000000100: n5504 = n5502;
      13'b0000000000010: n5504 = n5497;
      13'b0000000000001: n5504 = n5502;
      default: n5504 = 1'bX;
    endcase
  assign n5505 = n2762[27]; // extract
  assign n5506 = n4028[27]; // extract
  assign n5507 = n5072[27]; // extract
  assign n5508 = n5318[27]; // extract
  assign n5509 = fpsr[27]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5511 = n5508;
      13'b0100000000000: n5511 = n5509;
      13'b0010000000000: n5511 = n5507;
      13'b0001000000000: n5511 = n5509;
      13'b0000100000000: n5511 = n5509;
      13'b0000010000000: n5511 = n5509;
      13'b0000001000000: n5511 = n5509;
      13'b0000000100000: n5511 = n5509;
      13'b0000000010000: n5511 = n5509;
      13'b0000000001000: n5511 = n5506;
      13'b0000000000100: n5511 = n5509;
      13'b0000000000010: n5511 = n5505;
      13'b0000000000001: n5511 = n5509;
      default: n5511 = 1'bX;
    endcase
  assign n5512 = n2762[31:28]; // extract
  assign n5513 = n4028[31:28]; // extract
  assign n5514 = n5072[31:28]; // extract
  assign n5515 = n5318[31:28]; // extract
  assign n5516 = fpsr[31:28]; // extract
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5518 = n5515;
      13'b0100000000000: n5518 = n5516;
      13'b0010000000000: n5518 = n5514;
      13'b0001000000000: n5518 = n5516;
      13'b0000100000000: n5518 = n5516;
      13'b0000010000000: n5518 = n5516;
      13'b0000001000000: n5518 = n4342;
      13'b0000000100000: n5518 = n5516;
      13'b0000000010000: n5518 = n5516;
      13'b0000000001000: n5518 = n5513;
      13'b0000000000100: n5518 = n3628;
      13'b0000000000010: n5518 = n5512;
      13'b0000000000001: n5518 = n5516;
      default: n5518 = 4'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5522 = n5320;
      13'b0100000000000: n5522 = fpiar;
      13'b0010000000000: n5522 = n5074;
      13'b0001000000000: n5522 = fpiar;
      13'b0000100000000: n5522 = fpiar;
      13'b0000010000000: n5522 = fpiar;
      13'b0000001000000: n5522 = fpiar;
      13'b0000000100000: n5522 = fpiar;
      13'b0000000010000: n5522 = fpiar;
      13'b0000000001000: n5522 = fpiar;
      13'b0000000000100: n5522 = fpiar;
      13'b0000000000010: n5522 = n2763;
      13'b0000000000001: n5522 = fpiar;
      default: n5522 = 32'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5526 = n5322;
      13'b0100000000000: n5526 = fpcr_rounding_mode_valid;
      13'b0010000000000: n5526 = n5075;
      13'b0001000000000: n5526 = fpcr_rounding_mode_valid;
      13'b0000100000000: n5526 = fpcr_rounding_mode_valid;
      13'b0000010000000: n5526 = fpcr_rounding_mode_valid;
      13'b0000001000000: n5526 = fpcr_rounding_mode_valid;
      13'b0000000100000: n5526 = fpcr_rounding_mode_valid;
      13'b0000000010000: n5526 = fpcr_rounding_mode_valid;
      13'b0000000001000: n5526 = n3667;
      13'b0000000000100: n5526 = fpcr_rounding_mode_valid;
      13'b0000000000010: n5526 = fpcr_rounding_mode_valid;
      13'b0000000000001: n5526 = fpcr_rounding_mode_valid;
      default: n5526 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5528 = n5323;
      13'b0100000000000: n5528 = fpcr_precision_valid;
      13'b0010000000000: n5528 = n5076;
      13'b0001000000000: n5528 = fpcr_precision_valid;
      13'b0000100000000: n5528 = fpcr_precision_valid;
      13'b0000010000000: n5528 = fpcr_precision_valid;
      13'b0000001000000: n5528 = fpcr_precision_valid;
      13'b0000000100000: n5528 = fpcr_precision_valid;
      13'b0000000010000: n5528 = fpcr_precision_valid;
      13'b0000000001000: n5528 = n4029;
      13'b0000000000100: n5528 = fpcr_precision_valid;
      13'b0000000000010: n5528 = fpcr_precision_valid;
      13'b0000000000001: n5528 = fpcr_precision_valid;
      default: n5528 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5530 = fpcr_precision_bits;
      13'b0100000000000: n5530 = fpcr_precision_bits;
      13'b0010000000000: n5530 = fpcr_precision_bits;
      13'b0001000000000: n5530 = fpcr_precision_bits;
      13'b0000100000000: n5530 = fpcr_precision_bits;
      13'b0000010000000: n5530 = fpcr_precision_bits;
      13'b0000001000000: n5530 = fpcr_precision_bits;
      13'b0000000100000: n5530 = fpcr_precision_bits;
      13'b0000000010000: n5530 = fpcr_precision_bits;
      13'b0000000001000: n5530 = n4030;
      13'b0000000000100: n5530 = fpcr_precision_bits;
      13'b0000000000010: n5530 = fpcr_precision_bits;
      13'b0000000000001: n5530 = fpcr_precision_bits;
      default: n5530 = 2'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5534 = restore_privilege_violation;
      13'b0100000000000: n5534 = restore_privilege_violation;
      13'b0010000000000: n5534 = restore_privilege_violation;
      13'b0001000000000: n5534 = restore_privilege_violation;
      13'b0000100000000: n5534 = restore_privilege_violation;
      13'b0000010000000: n5534 = restore_privilege_violation;
      13'b0000001000000: n5534 = restore_privilege_violation;
      13'b0000000100000: n5534 = restore_privilege_violation;
      13'b0000000010000: n5534 = restore_privilege_violation;
      13'b0000000001000: n5534 = restore_privilege_violation;
      13'b0000000000100: n5534 = restore_privilege_violation;
      13'b0000000000010: n5534 = n911;
      13'b0000000000001: n5534 = restore_privilege_violation;
      default: n5534 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5536 = operation_word_cir;
      13'b0100000000000: n5536 = operation_word_cir;
      13'b0010000000000: n5536 = operation_word_cir;
      13'b0001000000000: n5536 = operation_word_cir;
      13'b0000100000000: n5536 = operation_word_cir;
      13'b0000010000000: n5536 = operation_word_cir;
      13'b0000001000000: n5536 = operation_word_cir;
      13'b0000000100000: n5536 = operation_word_cir;
      13'b0000000010000: n5536 = operation_word_cir;
      13'b0000000001000: n5536 = operation_word_cir;
      13'b0000000000100: n5536 = operation_word_cir;
      13'b0000000000010: n5536 = n2764;
      13'b0000000000001: n5536 = operation_word_cir;
      default: n5536 = 16'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5538 = command_address_cir;
      13'b0100000000000: n5538 = command_address_cir;
      13'b0010000000000: n5538 = command_address_cir;
      13'b0001000000000: n5538 = command_address_cir;
      13'b0000100000000: n5538 = command_address_cir;
      13'b0000010000000: n5538 = command_address_cir;
      13'b0000001000000: n5538 = command_address_cir;
      13'b0000000100000: n5538 = command_address_cir;
      13'b0000000010000: n5538 = command_address_cir;
      13'b0000000001000: n5538 = command_address_cir;
      13'b0000000000100: n5538 = command_address_cir;
      13'b0000000000010: n5538 = n2765;
      13'b0000000000001: n5538 = command_address_cir;
      default: n5538 = 32'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5544 = n5330;
      13'b0100000000000: n5544 = n5176;
      13'b0010000000000: n5544 = n5078;
      13'b0001000000000: n5544 = n4588;
      13'b0000100000000: n5544 = 4'b0000;
      13'b0000010000000: n5544 = 4'b0000;
      13'b0000001000000: n5544 = n4344;
      13'b0000000100000: n5544 = 4'b0000;
      13'b0000000010000: n5544 = 4'b0000;
      13'b0000000001000: n5544 = n4032;
      13'b0000000000100: n5544 = n3630;
      13'b0000000000010: n5544 = n2766;
      13'b0000000000001: n5544 = n846;
      default: n5544 = 4'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5548 = fsave_frame_format_latched;
      13'b0100000000000: n5548 = fsave_frame_format_latched;
      13'b0010000000000: n5548 = fsave_frame_format_latched;
      13'b0001000000000: n5548 = fsave_frame_format_latched;
      13'b0000100000000: n5548 = fsave_frame_format_latched;
      13'b0000010000000: n5548 = fsave_frame_format_latched;
      13'b0000001000000: n5548 = fsave_frame_format_latched;
      13'b0000000100000: n5548 = fsave_frame_format_latched;
      13'b0000000010000: n5548 = fsave_frame_format_latched;
      13'b0000000001000: n5548 = fsave_frame_format_latched;
      13'b0000000000100: n5548 = fsave_frame_format_latched;
      13'b0000000000010: n5548 = n2768;
      13'b0000000000001: n5548 = n848;
      default: n5548 = 8'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5551 = fpu_just_reset;
      13'b0100000000000: n5551 = fpu_just_reset;
      13'b0010000000000: n5551 = n5079;
      13'b0001000000000: n5551 = fpu_just_reset;
      13'b0000100000000: n5551 = fpu_just_reset;
      13'b0000010000000: n5551 = fpu_just_reset;
      13'b0000001000000: n5551 = fpu_just_reset;
      13'b0000000100000: n5551 = fpu_just_reset;
      13'b0000000010000: n5551 = fpu_just_reset;
      13'b0000000001000: n5551 = fpu_just_reset;
      13'b0000000000100: n5551 = fpu_just_reset;
      13'b0000000000010: n5551 = 1'b0;
      13'b0000000000001: n5551 = fpu_just_reset;
      default: n5551 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5553 = movem_register_list;
      13'b0100000000000: n5553 = movem_register_list;
      13'b0010000000000: n5553 = movem_register_list;
      13'b0001000000000: n5553 = movem_register_list;
      13'b0000100000000: n5553 = movem_register_list;
      13'b0000010000000: n5553 = movem_register_list;
      13'b0000001000000: n5553 = movem_register_list;
      13'b0000000100000: n5553 = movem_register_list;
      13'b0000000010000: n5553 = movem_register_list;
      13'b0000000001000: n5553 = movem_register_list;
      13'b0000000000100: n5553 = movem_register_list;
      13'b0000000000010: n5553 = n2769;
      13'b0000000000001: n5553 = movem_register_list;
      default: n5553 = 8'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5555 = movem_direction;
      13'b0100000000000: n5555 = movem_direction;
      13'b0010000000000: n5555 = movem_direction;
      13'b0001000000000: n5555 = movem_direction;
      13'b0000100000000: n5555 = movem_direction;
      13'b0000010000000: n5555 = movem_direction;
      13'b0000001000000: n5555 = movem_direction;
      13'b0000000100000: n5555 = movem_direction;
      13'b0000000010000: n5555 = movem_direction;
      13'b0000000001000: n5555 = movem_direction;
      13'b0000000000100: n5555 = movem_direction;
      13'b0000000000010: n5555 = n2770;
      13'b0000000000001: n5555 = movem_direction;
      default: n5555 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5559 = timeout_counter;
      13'b0100000000000: n5559 = timeout_counter;
      13'b0010000000000: n5559 = timeout_counter;
      13'b0001000000000: n5559 = timeout_counter;
      13'b0000100000000: n5559 = timeout_counter;
      13'b0000010000000: n5559 = timeout_counter;
      13'b0000001000000: n5559 = timeout_counter;
      13'b0000000100000: n5559 = timeout_counter;
      13'b0000000010000: n5559 = timeout_counter;
      13'b0000000001000: n5559 = n4034;
      13'b0000000000100: n5559 = 8'b00000000;
      13'b0000000000010: n5559 = 8'b00000000;
      13'b0000000000001: n5559 = timeout_counter;
      default: n5559 = 8'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5561 = fsave_counter;
      13'b0100000000000: n5561 = fsave_counter;
      13'b0010000000000: n5561 = n5080;
      13'b0001000000000: n5561 = fsave_counter;
      13'b0000100000000: n5561 = fsave_counter;
      13'b0000010000000: n5561 = fsave_counter;
      13'b0000001000000: n5561 = fsave_counter;
      13'b0000000100000: n5561 = fsave_counter;
      13'b0000000010000: n5561 = fsave_counter;
      13'b0000000001000: n5561 = fsave_counter;
      13'b0000000000100: n5561 = fsave_counter;
      13'b0000000000010: n5561 = n2771;
      13'b0000000000001: n5561 = n849;
      default: n5561 = 6'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5563 = frestore_frame_format;
      13'b0100000000000: n5563 = frestore_frame_format;
      13'b0010000000000: n5563 = n5081;
      13'b0001000000000: n5563 = frestore_frame_format;
      13'b0000100000000: n5563 = frestore_frame_format;
      13'b0000010000000: n5563 = frestore_frame_format;
      13'b0000001000000: n5563 = frestore_frame_format;
      13'b0000000100000: n5563 = frestore_frame_format;
      13'b0000000010000: n5563 = frestore_frame_format;
      13'b0000000001000: n5563 = frestore_frame_format;
      13'b0000000000100: n5563 = frestore_frame_format;
      13'b0000000000010: n5563 = n2772;
      13'b0000000000001: n5563 = n850;
      default: n5563 = 8'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5569 = frestore_fp_temp;
      13'b0100000000000: n5569 = frestore_fp_temp;
      13'b0010000000000: n5569 = n5082;
      13'b0001000000000: n5569 = frestore_fp_temp;
      13'b0000100000000: n5569 = frestore_fp_temp;
      13'b0000010000000: n5569 = frestore_fp_temp;
      13'b0000001000000: n5569 = frestore_fp_temp;
      13'b0000000100000: n5569 = frestore_fp_temp;
      13'b0000000010000: n5569 = frestore_fp_temp;
      13'b0000000001000: n5569 = frestore_fp_temp;
      13'b0000000000100: n5569 = frestore_fp_temp;
      13'b0000000000010: n5569 = frestore_fp_temp;
      13'b0000000000001: n5569 = frestore_fp_temp;
      default: n5569 = 640'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5571 = exception_code_internal;
      13'b0100000000000: n5571 = exception_code_internal;
      13'b0010000000000: n5571 = n5083;
      13'b0001000000000: n5571 = exception_code_internal;
      13'b0000100000000: n5571 = exception_code_internal;
      13'b0000010000000: n5571 = exception_code_internal;
      13'b0000001000000: n5571 = n4075;
      13'b0000000100000: n5571 = exception_code_internal;
      13'b0000000010000: n5571 = exception_code_internal;
      13'b0000000001000: n5571 = n4035;
      13'b0000000000100: n5571 = n3631;
      13'b0000000000010: n5571 = n2775;
      13'b0000000000001: n5571 = n853;
      default: n5571 = 8'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5574 = alu_start_operation;
      13'b0100000000000: n5574 = alu_start_operation;
      13'b0010000000000: n5574 = alu_start_operation;
      13'b0001000000000: n5574 = alu_start_operation;
      13'b0000100000000: n5574 = alu_start_operation;
      13'b0000010000000: n5574 = alu_start_operation;
      13'b0000001000000: n5574 = alu_start_operation;
      13'b0000000100000: n5574 = alu_start_operation;
      13'b0000000010000: n5574 = alu_start_operation;
      13'b0000000001000: n5574 = 1'b0;
      13'b0000000000100: n5574 = n3633;
      13'b0000000000010: n5574 = alu_start_operation;
      13'b0000000000001: n5574 = alu_start_operation;
      default: n5574 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5576 = alu_operation_code;
      13'b0100000000000: n5576 = alu_operation_code;
      13'b0010000000000: n5576 = alu_operation_code;
      13'b0001000000000: n5576 = alu_operation_code;
      13'b0000100000000: n5576 = alu_operation_code;
      13'b0000010000000: n5576 = alu_operation_code;
      13'b0000001000000: n5576 = alu_operation_code;
      13'b0000000100000: n5576 = alu_operation_code;
      13'b0000000010000: n5576 = alu_operation_code;
      13'b0000000001000: n5576 = alu_operation_code;
      13'b0000000000100: n5576 = n3635;
      13'b0000000000010: n5576 = alu_operation_code;
      13'b0000000000001: n5576 = alu_operation_code;
      default: n5576 = 7'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5578 = alu_operand_a;
      13'b0100000000000: n5578 = alu_operand_a;
      13'b0010000000000: n5578 = alu_operand_a;
      13'b0001000000000: n5578 = alu_operand_a;
      13'b0000100000000: n5578 = alu_operand_a;
      13'b0000010000000: n5578 = alu_operand_a;
      13'b0000001000000: n5578 = alu_operand_a;
      13'b0000000100000: n5578 = alu_operand_a;
      13'b0000000010000: n5578 = alu_operand_a;
      13'b0000000001000: n5578 = alu_operand_a;
      13'b0000000000100: n5578 = n3636;
      13'b0000000000010: n5578 = alu_operand_a;
      13'b0000000000001: n5578 = alu_operand_a;
      default: n5578 = 80'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5580 = alu_operand_b;
      13'b0100000000000: n5580 = alu_operand_b;
      13'b0010000000000: n5580 = alu_operand_b;
      13'b0001000000000: n5580 = alu_operand_b;
      13'b0000100000000: n5580 = alu_operand_b;
      13'b0000010000000: n5580 = alu_operand_b;
      13'b0000001000000: n5580 = alu_operand_b;
      13'b0000000100000: n5580 = alu_operand_b;
      13'b0000000010000: n5580 = alu_operand_b;
      13'b0000000001000: n5580 = alu_operand_b;
      13'b0000000000100: n5580 = n3637;
      13'b0000000000010: n5580 = alu_operand_b;
      13'b0000000000001: n5580 = alu_operand_b;
      default: n5580 = 80'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5583 = trans_start_operation;
      13'b0100000000000: n5583 = trans_start_operation;
      13'b0010000000000: n5583 = trans_start_operation;
      13'b0001000000000: n5583 = trans_start_operation;
      13'b0000100000000: n5583 = trans_start_operation;
      13'b0000010000000: n5583 = trans_start_operation;
      13'b0000001000000: n5583 = trans_start_operation;
      13'b0000000100000: n5583 = trans_start_operation;
      13'b0000000010000: n5583 = trans_start_operation;
      13'b0000000001000: n5583 = 1'b0;
      13'b0000000000100: n5583 = n3638;
      13'b0000000000010: n5583 = trans_start_operation;
      13'b0000000000001: n5583 = trans_start_operation;
      default: n5583 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5585 = trans_operation_code;
      13'b0100000000000: n5585 = trans_operation_code;
      13'b0010000000000: n5585 = trans_operation_code;
      13'b0001000000000: n5585 = trans_operation_code;
      13'b0000100000000: n5585 = trans_operation_code;
      13'b0000010000000: n5585 = trans_operation_code;
      13'b0000001000000: n5585 = trans_operation_code;
      13'b0000000100000: n5585 = trans_operation_code;
      13'b0000000010000: n5585 = trans_operation_code;
      13'b0000000001000: n5585 = trans_operation_code;
      13'b0000000000100: n5585 = n3639;
      13'b0000000000010: n5585 = trans_operation_code;
      13'b0000000000001: n5585 = trans_operation_code;
      default: n5585 = 7'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5587 = trans_operand;
      13'b0100000000000: n5587 = trans_operand;
      13'b0010000000000: n5587 = trans_operand;
      13'b0001000000000: n5587 = trans_operand;
      13'b0000100000000: n5587 = trans_operand;
      13'b0000010000000: n5587 = trans_operand;
      13'b0000001000000: n5587 = trans_operand;
      13'b0000000100000: n5587 = trans_operand;
      13'b0000000010000: n5587 = trans_operand;
      13'b0000000001000: n5587 = trans_operand;
      13'b0000000000100: n5587 = n3640;
      13'b0000000000010: n5587 = trans_operand;
      13'b0000000000001: n5587 = trans_operand;
      default: n5587 = 80'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5589 = final_result;
      13'b0100000000000: n5589 = final_result;
      13'b0010000000000: n5589 = final_result;
      13'b0001000000000: n5589 = final_result;
      13'b0000100000000: n5589 = final_result;
      13'b0000010000000: n5589 = final_result;
      13'b0000001000000: n5589 = final_result;
      13'b0000000100000: n5589 = final_result;
      13'b0000000010000: n5589 = final_result;
      13'b0000000001000: n5589 = n4036;
      13'b0000000000100: n5589 = final_result;
      13'b0000000000010: n5589 = final_result;
      13'b0000000000001: n5589 = final_result;
      default: n5589 = 80'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5591 = final_overflow;
      13'b0100000000000: n5591 = final_overflow;
      13'b0010000000000: n5591 = final_overflow;
      13'b0001000000000: n5591 = final_overflow;
      13'b0000100000000: n5591 = final_overflow;
      13'b0000010000000: n5591 = final_overflow;
      13'b0000001000000: n5591 = final_overflow;
      13'b0000000100000: n5591 = final_overflow;
      13'b0000000010000: n5591 = final_overflow;
      13'b0000000001000: n5591 = n4037;
      13'b0000000000100: n5591 = final_overflow;
      13'b0000000000010: n5591 = final_overflow;
      13'b0000000000001: n5591 = final_overflow;
      default: n5591 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5593 = final_underflow;
      13'b0100000000000: n5593 = final_underflow;
      13'b0010000000000: n5593 = final_underflow;
      13'b0001000000000: n5593 = final_underflow;
      13'b0000100000000: n5593 = final_underflow;
      13'b0000010000000: n5593 = final_underflow;
      13'b0000001000000: n5593 = final_underflow;
      13'b0000000100000: n5593 = final_underflow;
      13'b0000000010000: n5593 = final_underflow;
      13'b0000000001000: n5593 = n4038;
      13'b0000000000100: n5593 = final_underflow;
      13'b0000000000010: n5593 = final_underflow;
      13'b0000000000001: n5593 = final_underflow;
      default: n5593 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5595 = final_inexact;
      13'b0100000000000: n5595 = final_inexact;
      13'b0010000000000: n5595 = final_inexact;
      13'b0001000000000: n5595 = final_inexact;
      13'b0000100000000: n5595 = final_inexact;
      13'b0000010000000: n5595 = final_inexact;
      13'b0000001000000: n5595 = final_inexact;
      13'b0000000100000: n5595 = final_inexact;
      13'b0000000010000: n5595 = final_inexact;
      13'b0000000001000: n5595 = n4039;
      13'b0000000000100: n5595 = final_inexact;
      13'b0000000000010: n5595 = final_inexact;
      13'b0000000000001: n5595 = final_inexact;
      default: n5595 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5597 = final_invalid;
      13'b0100000000000: n5597 = final_invalid;
      13'b0010000000000: n5597 = final_invalid;
      13'b0001000000000: n5597 = final_invalid;
      13'b0000100000000: n5597 = final_invalid;
      13'b0000010000000: n5597 = final_invalid;
      13'b0000001000000: n5597 = final_invalid;
      13'b0000000100000: n5597 = final_invalid;
      13'b0000000010000: n5597 = final_invalid;
      13'b0000000001000: n5597 = n4040;
      13'b0000000000100: n5597 = final_invalid;
      13'b0000000000010: n5597 = final_invalid;
      13'b0000000000001: n5597 = final_invalid;
      default: n5597 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5599 = result_data;
      13'b0100000000000: n5599 = result_data;
      13'b0010000000000: n5599 = result_data;
      13'b0001000000000: n5599 = result_data;
      13'b0000100000000: n5599 = result_data;
      13'b0000010000000: n5599 = result_data;
      13'b0000001000000: n5599 = result_data;
      13'b0000000100000: n5599 = result_data;
      13'b0000000010000: n5599 = result_data;
      13'b0000000001000: n5599 = n4041;
      13'b0000000000100: n5599 = n3641;
      13'b0000000000010: n5599 = result_data;
      13'b0000000000001: n5599 = result_data;
      default: n5599 = 80'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5601 = converter_start;
      13'b0100000000000: n5601 = converter_start;
      13'b0010000000000: n5601 = converter_start;
      13'b0001000000000: n5601 = converter_start;
      13'b0000100000000: n5601 = converter_start;
      13'b0000010000000: n5601 = converter_start;
      13'b0000001000000: n5601 = converter_start;
      13'b0000000100000: n5601 = converter_start;
      13'b0000000010000: n5601 = converter_start;
      13'b0000000001000: n5601 = converter_start;
      13'b0000000000100: n5601 = converter_start;
      13'b0000000000010: n5601 = n2776;
      13'b0000000000001: n5601 = converter_start;
      default: n5601 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5603 = converter_source_format;
      13'b0100000000000: n5603 = converter_source_format;
      13'b0010000000000: n5603 = converter_source_format;
      13'b0001000000000: n5603 = converter_source_format;
      13'b0000100000000: n5603 = converter_source_format;
      13'b0000010000000: n5603 = converter_source_format;
      13'b0000001000000: n5603 = converter_source_format;
      13'b0000000100000: n5603 = converter_source_format;
      13'b0000000010000: n5603 = converter_source_format;
      13'b0000000001000: n5603 = converter_source_format;
      13'b0000000000100: n5603 = converter_source_format;
      13'b0000000000010: n5603 = n2777;
      13'b0000000000001: n5603 = converter_source_format;
      default: n5603 = 3'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5605 = converter_dest_format;
      13'b0100000000000: n5605 = converter_dest_format;
      13'b0010000000000: n5605 = converter_dest_format;
      13'b0001000000000: n5605 = converter_dest_format;
      13'b0000100000000: n5605 = converter_dest_format;
      13'b0000010000000: n5605 = converter_dest_format;
      13'b0000001000000: n5605 = converter_dest_format;
      13'b0000000100000: n5605 = converter_dest_format;
      13'b0000000010000: n5605 = converter_dest_format;
      13'b0000000001000: n5605 = converter_dest_format;
      13'b0000000000100: n5605 = converter_dest_format;
      13'b0000000000010: n5605 = n2778;
      13'b0000000000001: n5605 = converter_dest_format;
      default: n5605 = 3'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5607 = converter_data_in;
      13'b0100000000000: n5607 = converter_data_in;
      13'b0010000000000: n5607 = converter_data_in;
      13'b0001000000000: n5607 = converter_data_in;
      13'b0000100000000: n5607 = converter_data_in;
      13'b0000010000000: n5607 = converter_data_in;
      13'b0000001000000: n5607 = converter_data_in;
      13'b0000000100000: n5607 = converter_data_in;
      13'b0000000010000: n5607 = converter_data_in;
      13'b0000000001000: n5607 = converter_data_in;
      13'b0000000000100: n5607 = converter_data_in;
      13'b0000000000010: n5607 = n2779;
      13'b0000000000001: n5607 = converter_data_in;
      default: n5607 = 96'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5609 = rom_offset;
      13'b0100000000000: n5609 = rom_offset;
      13'b0010000000000: n5609 = rom_offset;
      13'b0001000000000: n5609 = rom_offset;
      13'b0000100000000: n5609 = rom_offset;
      13'b0000010000000: n5609 = rom_offset;
      13'b0000001000000: n5609 = rom_offset;
      13'b0000000100000: n5609 = rom_offset;
      13'b0000000010000: n5609 = rom_offset;
      13'b0000000001000: n5609 = rom_offset;
      13'b0000000000100: n5609 = rom_offset;
      13'b0000000000010: n5609 = n2780;
      13'b0000000000001: n5609 = rom_offset;
      default: n5609 = 7'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5611 = rom_read_enable;
      13'b0100000000000: n5611 = rom_read_enable;
      13'b0010000000000: n5611 = rom_read_enable;
      13'b0001000000000: n5611 = rom_read_enable;
      13'b0000100000000: n5611 = rom_read_enable;
      13'b0000010000000: n5611 = rom_read_enable;
      13'b0000001000000: n5611 = n4077;
      13'b0000000100000: n5611 = rom_read_enable;
      13'b0000000010000: n5611 = rom_read_enable;
      13'b0000000001000: n5611 = rom_read_enable;
      13'b0000000000100: n5611 = rom_read_enable;
      13'b0000000000010: n5611 = n2781;
      13'b0000000000001: n5611 = rom_read_enable;
      default: n5611 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5613 = movem_predecrement;
      13'b0100000000000: n5613 = movem_predecrement;
      13'b0010000000000: n5613 = movem_predecrement;
      13'b0001000000000: n5613 = movem_predecrement;
      13'b0000100000000: n5613 = movem_predecrement;
      13'b0000010000000: n5613 = movem_predecrement;
      13'b0000001000000: n5613 = movem_predecrement;
      13'b0000000100000: n5613 = movem_predecrement;
      13'b0000000010000: n5613 = movem_predecrement;
      13'b0000000001000: n5613 = movem_predecrement;
      13'b0000000000100: n5613 = movem_predecrement;
      13'b0000000000010: n5613 = n2782;
      13'b0000000000001: n5613 = movem_predecrement;
      default: n5613 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5615 = movem_postincrement;
      13'b0100000000000: n5615 = movem_postincrement;
      13'b0010000000000: n5615 = movem_postincrement;
      13'b0001000000000: n5615 = movem_postincrement;
      13'b0000100000000: n5615 = movem_postincrement;
      13'b0000010000000: n5615 = movem_postincrement;
      13'b0000001000000: n5615 = movem_postincrement;
      13'b0000000100000: n5615 = movem_postincrement;
      13'b0000000010000: n5615 = movem_postincrement;
      13'b0000000001000: n5615 = movem_postincrement;
      13'b0000000000100: n5615 = movem_postincrement;
      13'b0000000000010: n5615 = n2783;
      13'b0000000000001: n5615 = movem_postincrement;
      default: n5615 = 1'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5623 = fp_to_int_shift;
      13'b0100000000000: n5623 = fp_to_int_shift;
      13'b0010000000000: n5623 = fp_to_int_shift;
      13'b0001000000000: n5623 = fp_to_int_shift;
      13'b0000100000000: n5623 = fp_to_int_shift;
      13'b0000010000000: n5623 = fp_to_int_shift;
      13'b0000001000000: n5623 = fp_to_int_shift;
      13'b0000000100000: n5623 = fp_to_int_shift;
      13'b0000000010000: n5623 = fp_to_int_shift;
      13'b0000000001000: n5623 = fp_to_int_shift;
      13'b0000000000100: n5623 = fp_to_int_shift;
      13'b0000000000010: n5623 = n2787;
      13'b0000000000001: n5623 = fp_to_int_shift;
      default: n5623 = 6'bX;
    endcase
  /* TG68K_FPU.vhd:1240:33  */
  always @*
    case (n5333)
      13'b1000000000000: n5625 = fp_to_int_result;
      13'b0100000000000: n5625 = fp_to_int_result;
      13'b0010000000000: n5625 = fp_to_int_result;
      13'b0001000000000: n5625 = fp_to_int_result;
      13'b0000100000000: n5625 = fp_to_int_result;
      13'b0000010000000: n5625 = fp_to_int_result;
      13'b0000001000000: n5625 = fp_to_int_result;
      13'b0000000100000: n5625 = fp_to_int_result;
      13'b0000000010000: n5625 = fp_to_int_result;
      13'b0000000001000: n5625 = fp_to_int_result;
      13'b0000000000100: n5625 = fp_to_int_result;
      13'b0000000000010: n5625 = n2788;
      13'b0000000000001: n5625 = fp_to_int_result;
      default: n5625 = 32'bX;
    endcase
  /* TG68K_FPU.vhd:3507:52  */
  assign n5626 = cir_read | cir_write;
  /* TG68K_FPU.vhd:3507:76  */
  assign n5627 = {26'b0, cir_address};  //  uext
  /* TG68K_FPU.vhd:3507:110  */
  assign n5628 = {1'b0, n5627};  //  uext
  /* TG68K_FPU.vhd:3507:110  */
  assign n5630 = $signed(n5628) > $signed(32'b00000000000000000000000000001000);
  /* TG68K_FPU.vhd:3507:72  */
  assign n5631 = n5630 & n5626;
  /* TG68K_FPU.vhd:3507:33  */
  assign n5633 = n5631 ? 1'b1 : n5344;
  /* TG68K_FPU.vhd:3507:33  */
  assign n5635 = n5631 ? 8'b00001110 : n5571;
  /* TG68K_FPU.vhd:3516:49  */
  assign n5637 = cir_address == 5'b00000;
  /* TG68K_FPU.vhd:3519:49  */
  assign n5639 = cir_address == 5'b00010;
  /* TG68K_FPU.vhd:3522:49  */
  assign n5641 = cir_address == 5'b00011;
  /* TG68K_FPU.vhd:3525:49  */
  assign n5643 = cir_address == 5'b00110;
  /* TG68K_FPU.vhd:3528:49  */
  assign n5645 = cir_address == 5'b00111;
  /* TG68K_FPU.vhd:3528:62  */
  assign n5647 = cir_address == 5'b01000;
  /* TG68K_FPU.vhd:3528:62  */
  assign n5648 = n5645 | n5647;
  assign n5649 = {n5648, n5643, n5641, n5639, n5637};
  /* TG68K_FPU.vhd:3515:41  */
  always @*
    case (n5649)
      5'b10000: n5655 = 1'b1;
      5'b01000: n5655 = 1'b1;
      5'b00100: n5655 = 1'b1;
      5'b00010: n5655 = 1'b1;
      5'b00001: n5655 = 1'b1;
      default: n5655 = n5633;
    endcase
  /* TG68K_FPU.vhd:3515:41  */
  always @*
    case (n5649)
      5'b10000: n5661 = 8'b00001100;
      5'b01000: n5661 = 8'b00001100;
      5'b00100: n5661 = 8'b00001100;
      5'b00010: n5661 = 8'b00001100;
      5'b00001: n5661 = 8'b00001100;
      default: n5661 = n5635;
    endcase
  /* TG68K_FPU.vhd:3514:33  */
  assign n5662 = cir_write ? n5655 : n5633;
  /* TG68K_FPU.vhd:3514:33  */
  assign n5663 = cir_write ? n5661 : n5635;
  /* TG68K_FPU.vhd:3536:56  */
  assign n5664 = {29'b0, cir_handshake_state};  //  uext
  /* TG68K_FPU.vhd:3536:56  */
  assign n5666 = n5664 == 32'b00000000000000000000000000000110;
  /* TG68K_FPU.vhd:3542:41  */
  assign n5669 = cir_address_error ? 8'b00001110 : 8'b00001100;
  /* TG68K_FPU.vhd:3538:41  */
  assign n5671 = restore_privilege_violation ? 8'b00001000 : n5669;
  /* TG68K_FPU.vhd:3536:33  */
  assign n5673 = n5666 ? 1'b1 : n5662;
  /* TG68K_FPU.vhd:3536:33  */
  assign n5674 = n5666 ? n5671 : n5663;
  /* TG68K_FPU.vhd:3555:58  */
  assign n5675 = {22'b0, state_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3555:58  */
  assign n5677 = $signed(n5675) > $signed(32'b00000000000000000000001111101000);
  /* TG68K_FPU.vhd:3555:33  */
  assign n5679 = n5677 ? 1'b1 : n5673;
  /* TG68K_FPU.vhd:3555:33  */
  assign n5681 = n5677 ? 8'b00001111 : n5674;
  /* TG68K_FPU.vhd:3563:48  */
  assign n5683 = command_cir == 16'b0000000000000010;
  /* TG68K_FPU.vhd:3569:51  */
  assign n5685 = command_cir == 16'b0000000000000011;
  /* TG68K_FPU.vhd:3569:33  */
  assign n5687 = n5685 ? 1'b1 : n5342;
  /* TG68K_FPU.vhd:3569:33  */
  assign n5689 = n5685 ? 1'b0 : cir_address_error;
  /* TG68K_FPU.vhd:3569:33  */
  assign n5691 = n5685 ? 4'b0000 : n5544;
  /* TG68K_FPU.vhd:3563:33  */
  assign n5693 = n5683 ? 1'b0 : n5687;
  /* TG68K_FPU.vhd:3563:33  */
  assign n5695 = n5683 ? 1'b0 : n5679;
  /* TG68K_FPU.vhd:3563:33  */
  assign n5697 = n5683 ? 1'b0 : n5689;
  /* TG68K_FPU.vhd:3563:33  */
  assign n5699 = n5683 ? 4'b0000 : n5691;
  assign n5711 = {n5390, n5384, n5378, n5372, n5366};
  assign n5715 = {n5518, n5511, n5504, n5496, n5488, n5480, n5472, n5464, n5456, n5448, n5440, n5432, n5424, n5416, n5408, n5401};
  /* TG68K_FPU.vhd:3582:27  */
  assign n5934 = ~nReset;
  /* TG68K_FPU.vhd:3588:54  */
  assign n5937 = $unsigned(movem_reg_address) <= $unsigned(3'b111);
  /* TG68K_FPU.vhd:3589:75  */
  assign n5940 = 3'b111 - movem_reg_address;
  /* TG68K_FPU.vhd:3588:33  */
  assign n5944 = n5937 ? n7102 : 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* TG68K_FPU.vhd:3617:27  */
  assign n5953 = ~nReset;
  /* TG68K_FPU.vhd:3622:41  */
  assign n5956 = fpu_state == 4'b0000;
  /* TG68K_FPU.vhd:3621:33  */
  always @*
    case (n5956)
      1'b1: n5959 = 1'b0;
      default: n5959 = 1'b1;
    endcase
  /* TG68K_FPU.vhd:3635:27  */
  assign n5967 = ~nReset;
  /* TG68K_FPU.vhd:3671:33  */
  assign n5971 = supervisor_mode ? 3'b000 : 3'b011;
  /* TG68K_FPU.vhd:3687:68  */
  assign n5980 = ~cir_read_reg;
  /* TG68K_FPU.vhd:3687:51  */
  assign n5981 = n5980 & cir_read;
  /* TG68K_FPU.vhd:3690:48  */
  assign n5982 = ~cir_read;
  /* TG68K_FPU.vhd:3690:54  */
  assign n5983 = cir_read_reg & n5982;
  /* TG68K_FPU.vhd:3690:33  */
  assign n5987 = n5983 ? 1'b0 : cir_read_active;
  /* TG68K_FPU.vhd:3687:33  */
  assign n5991 = n5981 ? 1'b1 : n5987;
  /* TG68K_FPU.vhd:3696:58  */
  assign n5992 = cir_read_active | cir_write;
  /* TG68K_FPU.vhd:3697:84  */
  assign n5993 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3697:84  */
  assign n5995 = n5993 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3697:64  */
  assign n5996 = n5995[9:0];  // trunc
  /* TG68K_FPU.vhd:3699:64  */
  assign n5997 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3699:64  */
  assign n5999 = $signed(n5997) > $signed(32'b00000000000000000000001111101000);
  /* TG68K_FPU.vhd:3696:33  */
  assign n6005 = n6010 ? 1'b0 : n5991;
  /* TG68K_FPU.vhd:3699:41  */
  assign n6007 = n5999 ? 10'b0000000000 : n5996;
  /* TG68K_FPU.vhd:3696:33  */
  assign n6010 = n5999 & n5992;
  /* TG68K_FPU.vhd:3696:33  */
  assign n6012 = n5992 ? n6007 : 10'b0000000000;
  /* TG68K_FPU.vhd:3710:70  */
  assign n6013 = ~cir_write_reg;
  /* TG68K_FPU.vhd:3710:52  */
  assign n6014 = n6013 & cir_write;
  /* TG68K_FPU.vhd:3712:49  */
  assign n6026 = cir_address == 5'b00001;
  /* TG68K_FPU.vhd:3736:49  */
  assign n6048 = cir_address == 5'b00100;
  /* TG68K_FPU.vhd:3757:49  */
  assign n6081 = cir_address == 5'b00101;
  assign n6082 = {n6081, n6048, n6026};
  /* TG68K_FPU.vhd:3711:41  */
  always @*
    case (n6082)
      3'b100: n6083 = command_cir;
      3'b010: n6083 = command_cir;
      3'b001: n6083 = cir_data_in;
      default: n6083 = command_cir;
    endcase
  /* TG68K_FPU.vhd:3711:41  */
  always @*
    case (n6082)
      3'b100: n6087 = command_pending;
      3'b010: n6087 = command_pending;
      3'b001: n6087 = 1'b1;
      default: n6087 = command_pending;
    endcase
  /* TG68K_FPU.vhd:3710:33  */
  assign n6096 = n6014 ? n6087 : command_pending;
  /* TG68K_FPU.vhd:3787:33  */
  assign n6103 = cir_read ? 1'b1 : 1'b0;
  /* TG68K_FPU.vhd:3799:73  */
  assign n6105 = fpu_state == 4'b0001;
  /* TG68K_FPU.vhd:3799:99  */
  assign n6107 = fpu_state == 4'b1000;
  /* TG68K_FPU.vhd:3799:86  */
  assign n6108 = n6105 | n6107;
  /* TG68K_FPU.vhd:3799:121  */
  assign n6109 = n6108 | fpu_done_i;
  /* TG68K_FPU.vhd:3799:58  */
  assign n6110 = n6109 & command_pending;
  /* TG68K_FPU.vhd:3799:33  */
  assign n6112 = n6110 ? 1'b0 : n6096;
  /* TG68K_FPU.vhd:3813:67  */
  assign n6113 = cir_read | cir_write;
  /* TG68K_FPU.vhd:3813:49  */
  assign n6115 = n6113 ? 3'b001 : cir_handshake_state;
  /* TG68K_FPU.vhd:3806:41  */
  assign n6117 = cir_handshake_state == 3'b000;
  /* TG68K_FPU.vhd:3819:92  */
  assign n6118 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3819:92  */
  assign n6120 = n6118 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3819:72  */
  assign n6121 = n6120[9:0];  // trunc
  /* TG68K_FPU.vhd:3822:52  */
  assign n6122 = {26'b0, cir_address};  //  uext
  /* TG68K_FPU.vhd:3822:86  */
  assign n6123 = {1'b0, n6122};  //  uext
  /* TG68K_FPU.vhd:3822:86  */
  assign n6125 = $signed(n6123) > $signed(32'b00000000000000000000000000001000);
  /* TG68K_FPU.vhd:3826:68  */
  assign n6127 = cir_address == 5'b00011;
  /* TG68K_FPU.vhd:3826:93  */
  assign n6129 = cir_address == 5'b00100;
  /* TG68K_FPU.vhd:3826:78  */
  assign n6130 = n6127 | n6129;
  /* TG68K_FPU.vhd:3826:124  */
  assign n6131 = ~supervisor_mode;
  /* TG68K_FPU.vhd:3826:104  */
  assign n6132 = n6131 & n6130;
  /* TG68K_FPU.vhd:3832:88  */
  assign n6134 = cir_address == 5'b00000;
  /* TG68K_FPU.vhd:3832:113  */
  assign n6136 = cir_address == 5'b00001;
  /* TG68K_FPU.vhd:3832:98  */
  assign n6137 = n6134 | n6136;
  /* TG68K_FPU.vhd:3832:138  */
  assign n6139 = cir_address == 5'b00010;
  /* TG68K_FPU.vhd:3832:123  */
  assign n6140 = n6137 | n6139;
  /* TG68K_FPU.vhd:3832:71  */
  assign n6141 = n6140 & cir_write;
  /* TG68K_FPU.vhd:3832:49  */
  assign n6144 = n6141 ? 3'b110 : 3'b010;
  /* TG68K_FPU.vhd:3826:49  */
  assign n6148 = n6132 ? 3'b110 : n6144;
  /* TG68K_FPU.vhd:3822:49  */
  assign n6152 = n6125 ? 3'b110 : n6148;
  /* TG68K_FPU.vhd:3842:72  */
  assign n6155 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3842:72  */
  assign n6157 = $signed(n6155) > $signed(32'b00000000000000000000000001000000);
  /* TG68K_FPU.vhd:3842:49  */
  assign n6159 = n6157 ? 3'b110 : n6152;
  /* TG68K_FPU.vhd:3818:41  */
  assign n6163 = cir_handshake_state == 3'b001;
  /* TG68K_FPU.vhd:3848:92  */
  assign n6164 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3848:92  */
  assign n6166 = n6164 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3848:72  */
  assign n6167 = n6166[9:0];  // trunc
  /* TG68K_FPU.vhd:3855:49  */
  assign n6185 = cir_write ? 3'b011 : cir_handshake_state;
  /* TG68K_FPU.vhd:3850:49  */
  assign n6191 = cir_read ? 3'b011 : n6185;
  /* TG68K_FPU.vhd:3869:72  */
  assign n6196 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3869:72  */
  assign n6198 = $signed(n6196) > $signed(32'b00000000000000000000000010000000);
  /* TG68K_FPU.vhd:3869:49  */
  assign n6200 = n6198 ? 3'b110 : n6191;
  /* TG68K_FPU.vhd:3847:41  */
  assign n6204 = cir_handshake_state == 3'b010;
  /* TG68K_FPU.vhd:3874:41  */
  assign n6206 = cir_handshake_state == 3'b011;
  /* TG68K_FPU.vhd:3880:61  */
  assign n6207 = ~cir_read;
  /* TG68K_FPU.vhd:3880:81  */
  assign n6208 = ~cir_write;
  /* TG68K_FPU.vhd:3880:67  */
  assign n6209 = n6208 & n6207;
  /* TG68K_FPU.vhd:3880:49  */
  assign n6211 = n6209 ? 3'b101 : cir_handshake_state;
  /* TG68K_FPU.vhd:3885:72  */
  assign n6212 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3885:72  */
  assign n6214 = $signed(n6212) > $signed(32'b00000000000000000000000100000000);
  /* TG68K_FPU.vhd:3885:49  */
  assign n6216 = n6214 ? 3'b110 : n6211;
  /* TG68K_FPU.vhd:3878:41  */
  assign n6220 = cir_handshake_state == 3'b100;
  /* TG68K_FPU.vhd:3890:41  */
  assign n6222 = cir_handshake_state == 3'b101;
  /* TG68K_FPU.vhd:3909:72  */
  assign n6223 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3909:72  */
  assign n6225 = $signed(n6223) > $signed(32'b00000000000000000000000000100000);
  /* TG68K_FPU.vhd:3914:100  */
  assign n6226 = {22'b0, cir_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3914:100  */
  assign n6228 = n6226 + 32'b00000000000000000000000000000001;
  /* TG68K_FPU.vhd:3914:80  */
  assign n6229 = n6228[9:0];  // trunc
  /* TG68K_FPU.vhd:3909:49  */
  assign n6230 = n6225 ? n6012 : n6229;
  /* TG68K_FPU.vhd:3909:49  */
  assign n6232 = n6225 ? 3'b000 : cir_handshake_state;
  /* TG68K_FPU.vhd:3899:41  */
  assign n6238 = cir_handshake_state == 3'b110;
  assign n6239 = {n6238, n6222, n6220, n6206, n6204, n6163, n6117};
  /* TG68K_FPU.vhd:3805:33  */
  always @*
    case (n6239)
      7'b1000000: n6242 = n6230;
      7'b0100000: n6242 = 10'b0000000000;
      7'b0010000: n6242 = n6012;
      7'b0001000: n6242 = n6012;
      7'b0000100: n6242 = n6167;
      7'b0000010: n6242 = n6121;
      7'b0000001: n6242 = 10'b0000000000;
      default: n6242 = n6012;
    endcase
  /* TG68K_FPU.vhd:3805:33  */
  always @*
    case (n6239)
      7'b1000000: n6250 = n6232;
      7'b0100000: n6250 = 3'b000;
      7'b0010000: n6250 = n6216;
      7'b0001000: n6250 = 3'b100;
      7'b0000100: n6250 = n6200;
      7'b0000010: n6250 = n6159;
      7'b0000001: n6250 = n6115;
      default: n6250 = 3'b000;
    endcase
  /* TG68K_FPU.vhd:3925:41  */
  assign n6263 = fpu_state == 4'b0000;
  /* TG68K_FPU.vhd:3938:77  */
  assign n6265 = decoder_instruction_type == 4'b0000;
  /* TG68K_FPU.vhd:3943:81  */
  assign n6267 = decoder_source_format == 3'b110;
  /* TG68K_FPU.vhd:3943:98  */
  assign n6269 = decoder_source_format == 3'b100;
  /* TG68K_FPU.vhd:3943:98  */
  assign n6270 = n6267 | n6269;
  /* TG68K_FPU.vhd:3942:73  */
  always @*
    case (n6270)
      1'b1: n6273 = 16'b0000000000000001;
      default: n6273 = 16'b0000000000000000;
    endcase
  /* TG68K_FPU.vhd:3941:65  */
  assign n6275 = decoder_ea_mode == 3'b000;
  /* TG68K_FPU.vhd:3950:65  */
  assign n6277 = decoder_ea_mode == 3'b001;
  assign n6278 = {n6277, n6275};
  /* TG68K_FPU.vhd:3940:57  */
  always @*
    case (n6278)
      2'b10: n6281 = 16'b0000000000000001;
      2'b01: n6281 = n6273;
      default: n6281 = 16'b0000000000000000;
    endcase
  /* TG68K_FPU.vhd:3956:80  */
  assign n6283 = decoder_instruction_type == 4'b0001;
  /* TG68K_FPU.vhd:3959:80  */
  assign n6285 = decoder_instruction_type == 4'b0010;
  /* TG68K_FPU.vhd:3962:80  */
  assign n6287 = decoder_instruction_type == 4'b0100;
  /* TG68K_FPU.vhd:3964:76  */
  assign n6289 = decoder_ea_mode == 3'b000;
  /* TG68K_FPU.vhd:3964:57  */
  assign n6292 = n6289 ? 16'b0000000000000010 : 16'b0000000000000001;
  /* TG68K_FPU.vhd:3962:49  */
  assign n6294 = n6287 ? n6292 : 16'b0000000000000000;
  /* TG68K_FPU.vhd:3959:49  */
  assign n6296 = n6285 ? 16'b0000000000000001 : n6294;
  /* TG68K_FPU.vhd:3956:49  */
  assign n6298 = n6283 ? 16'b0000000000000010 : n6296;
  /* TG68K_FPU.vhd:3938:49  */
  assign n6299 = n6265 ? n6281 : n6298;
  /* TG68K_FPU.vhd:3936:41  */
  assign n6301 = fpu_state == 4'b0001;
  /* TG68K_FPU.vhd:3977:84  */
  assign n6303 = cir_address == 5'b00101;
  /* TG68K_FPU.vhd:3977:68  */
  assign n6304 = n6303 & cir_write;
  /* TG68K_FPU.vhd:3977:94  */
  assign n6305 = cir_data_valid_i & n6304;
  /* TG68K_FPU.vhd:3981:77  */
  assign n6306 = {22'b0, state_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:3981:77  */
  assign n6308 = $signed(n6306) > $signed(32'b00000000000000000000001111101000);
  /* TG68K_FPU.vhd:3981:49  */
  assign n6311 = n6308 ? 16'b0000000000000000 : 16'b0000000000000001;
  /* TG68K_FPU.vhd:3977:49  */
  assign n6313 = n6305 ? 16'b0000000000000000 : n6311;
  /* TG68K_FPU.vhd:3974:41  */
  assign n6315 = fpu_state == 4'b0010;
  /* TG68K_FPU.vhd:3991:41  */
  assign n6317 = fpu_state == 4'b0101;
  /* TG68K_FPU.vhd:3997:77  */
  assign n6319 = decoder_instruction_type == 4'b0001;
  /* TG68K_FPU.vhd:3999:91  */
  assign n6321 = cir_address == 5'b00110;
  /* TG68K_FPU.vhd:3999:75  */
  assign n6322 = n6321 & cir_read;
  /* TG68K_FPU.vhd:3999:101  */
  assign n6323 = cir_data_valid_i & n6322;
  /* TG68K_FPU.vhd:4003:85  */
  assign n6324 = {22'b0, state_timeout_counter};  //  uext
  /* TG68K_FPU.vhd:4003:85  */
  assign n6326 = $signed(n6324) > $signed(32'b00000000000000000000001111101000);
  /* TG68K_FPU.vhd:4003:57  */
  assign n6329 = n6326 ? 16'b0000000000000000 : 16'b0000000000000010;
  /* TG68K_FPU.vhd:3999:57  */
  assign n6331 = n6323 ? 16'b0000000000000000 : n6329;
  /* TG68K_FPU.vhd:3997:49  */
  assign n6333 = n6319 ? n6331 : 16'b0000000000000000;
  /* TG68K_FPU.vhd:3995:41  */
  assign n6335 = fpu_state == 4'b0110;
  /* TG68K_FPU.vhd:4018:41  */
  assign n6337 = fpu_state == 4'b0111;
  /* TG68K_FPU.vhd:4022:41  */
  assign n6339 = fpu_state == 4'b1000;
  assign n6343 = {n6339, n6337, n6335, n6317, n6315, n6301, n6263};
  /* TG68K_FPU.vhd:3924:33  */
  always @*
    case (n6343)
      7'b1000000: n6349 = 16'b0000000000000000;
      7'b0100000: n6349 = 16'b0000000000000000;
      7'b0010000: n6349 = n6333;
      7'b0001000: n6349 = 16'b0000000000000000;
      7'b0000100: n6349 = n6313;
      7'b0000010: n6349 = n6299;
      7'b0000001: n6349 = 16'b0000000000000000;
      default: n6349 = 16'b0000000000000000;
    endcase
  /* TG68K_FPU.vhd:4041:57  */
  assign n6350 = fpsr[31]; // extract
  assign n6352 = n6351[15:4]; // extract
  /* TG68K_FPU.vhd:4042:57  */
  assign n6354 = fpsr[30]; // extract
  /* TG68K_FPU.vhd:4043:57  */
  assign n6356 = fpsr[29]; // extract
  /* TG68K_FPU.vhd:4044:57  */
  assign n6358 = fpsr[28]; // extract
  /* TG68K_FPU.vhd:4050:46  */
  assign n6360 = fpu_state != 4'b0000;
  /* TG68K_FPU.vhd:4050:72  */
  assign n6362 = fpu_state != 4'b1001;
  /* TG68K_FPU.vhd:4050:58  */
  assign n6363 = n6362 & n6360;
  /* TG68K_FPU.vhd:4051:46  */
  assign n6365 = fpu_state != 4'b1010;
  /* TG68K_FPU.vhd:4050:91  */
  assign n6366 = n6365 & n6363;
  /* TG68K_FPU.vhd:4051:67  */
  assign n6367 = fpu_busy_internal & n6366;
  /* TG68K_FPU.vhd:4059:49  */
  assign n6369 = fsave_frame_format == 8'b00000000;
  /* TG68K_FPU.vhd:4060:49  */
  assign n6371 = fsave_frame_format == 8'b01100000;
  /* TG68K_FPU.vhd:4061:49  */
  assign n6373 = fsave_frame_format == 8'b11011000;
  assign n6374 = {n6373, n6371, n6369};
  /* TG68K_FPU.vhd:4058:41  */
  always @*
    case (n6374)
      3'b100: n6379 = 16'b1101100011010100;
      3'b010: n6379 = 16'b0110000000111000;
      3'b001: n6379 = 16'b0000000000000000;
      default: n6379 = 16'b0000000000000000;
    endcase
  /* TG68K_FPU.vhd:4050:33  */
  assign n6381 = n6367 ? 16'b0000000100000000 : n6379;
  /* TG68K_FPU.vhd:3664:25  */
  assign n6384 = n6014 & clkena;
  assign n6385 = {n6352, n6350, n6354, n6356, n6358};
  /* TG68K_FPU.vhd:4152:25  */
  assign n6530 = cir_address == 5'b00000;
  /* TG68K_FPU.vhd:4154:25  */
  assign n6532 = cir_address == 5'b00001;
  /* TG68K_FPU.vhd:4156:25  */
  assign n6534 = cir_address == 5'b00010;
  /* TG68K_FPU.vhd:4158:25  */
  assign n6536 = cir_address == 5'b00011;
  /* TG68K_FPU.vhd:4160:25  */
  assign n6538 = cir_address == 5'b00100;
  /* TG68K_FPU.vhd:4162:25  */
  assign n6540 = cir_address == 5'b00101;
  /* TG68K_FPU.vhd:4164:25  */
  assign n6542 = cir_address == 5'b00110;
  /* TG68K_FPU.vhd:4167:68  */
  assign n6543 = command_address_cir[15:0]; // extract
  /* TG68K_FPU.vhd:4166:25  */
  assign n6545 = cir_address == 5'b00111;
  /* TG68K_FPU.vhd:4169:68  */
  assign n6546 = command_address_cir[31:16]; // extract
  /* TG68K_FPU.vhd:4168:25  */
  assign n6548 = cir_address == 5'b01000;
  assign n6549 = {n6548, n6545, n6542, n6540, n6538, n6536, n6534, n6532, n6530};
  /* TG68K_FPU.vhd:4151:17  */
  always @*
    case (n6549)
      9'b100000000: n6554 = n6546;
      9'b010000000: n6554 = n6543;
      9'b001000000: n6554 = operation_word_cir;
      9'b000100000: n6554 = 16'bX;
      9'b000010000: n6554 = 16'bX;
      9'b000001000: n6554 = save_cir;
      9'b000000100: n6554 = condition_cir;
      9'b000000010: n6554 = 16'bX;
      9'b000000001: n6554 = response_cir;
      default: n6554 = 16'b0000000000000000;
    endcase
  /* TG68K_FPU.vhd:1230:17  */
  assign n6556 = clkena ? n5693 : fpu_done_i;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6557 <= 1'b0;
    else
      n6557 <= n6556;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6558 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6559 = clkena & n6558;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6560 = n6559 ? n5695 : fpu_exception_i;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6561 <= n6560;
  initial
    n6561 = 1'b0;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6562 = clkena ? n6103 : cir_data_valid_i;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6563 <= 1'b0;
    else
      n6563 <= n6562;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6564 = clkena ? n5346 : fp_registers;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6565 <= 640'b0111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000;
    else
      n6565 <= n6564;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6570 = clkena ? n5352 : fp_reg_write_enable;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6571 <= 1'b0;
    else
      n6571 <= n6570;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6572 = clkena ? n5354 : fp_reg_write_addr;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6573 <= 3'b000;
    else
      n6573 <= n6572;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6574 = clkena ? n5356 : fp_reg_write_data;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6575 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n6575 <= n6574;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6582 = clkena ? n5360 : fp_reg_access_valid;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6583 <= 1'b0;
    else
      n6583 <= n6582;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6588 = clkena ? n5711 : fpcr;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6589 <= 32'b00000000000000000000000000000000;
    else
      n6589 <= n6588;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6594 = clkena ? n5715 : fpsr;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6595 <= 32'b00000000000000000000000000000000;
    else
      n6595 <= n6594;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6598 = clkena ? n5522 : fpiar;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6599 <= 32'b00000000000000000000000000000000;
    else
      n6599 <= n6598;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6602 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6603 = clkena & n6602;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6604 = n6603 ? n5526 : fpcr_rounding_mode_valid;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6605 <= n6604;
  initial
    n6605 = 1'b1;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6606 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6607 = clkena & n6606;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6608 = n6607 ? n5528 : fpcr_precision_valid;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6609 <= n6608;
  initial
    n6609 = 1'b1;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6610 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6611 = clkena & n6610;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6612 = n6611 ? n5530 : fpcr_precision_bits;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6613 <= n6612;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6618 = clkena ? n6349 : response_cir;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6619 <= 16'b0000000000000000;
    else
      n6619 <= n6618;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6620 = n6384 ? n6083 : command_cir;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6621 <= 16'b0000000000000000;
    else
      n6621 <= n6620;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6622 = clkena ? n6385 : condition_cir;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6623 <= 16'b0000000000000000;
    else
      n6623 <= n6622;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6624 = clkena ? n6381 : save_cir;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6625 <= 16'b0000000000000000;
    else
      n6625 <= n6624;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6630 = clkena ? cir_read : cir_read_reg;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6631 <= 1'b0;
    else
      n6631 <= n6630;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6632 = clkena ? cir_write : cir_write_reg;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6633 <= 1'b0;
    else
      n6633 <= n6632;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6634 = clkena ? n6005 : cir_read_active;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6635 <= 1'b0;
    else
      n6635 <= n6634;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6636 = clkena ? n6242 : cir_timeout_counter;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6637 <= 10'b0000000000;
    else
      n6637 <= n6636;
  /* TG68K_FPU.vhd:1179:9  */
  always @(n743)
    n6638 <= 10'b0000000000;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6639 = clkena ? n6112 : command_pending;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6640 <= 1'b0;
    else
      n6640 <= n6639;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6643 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6644 = clkena & n6643;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6645 = n6644 ? n5534 : restore_privilege_violation;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6646 <= n6645;
  initial
    n6646 = 1'b0;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6653 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6654 = clkena & n6653;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6655 = n6654 ? n5697 : cir_address_error;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6656 <= n6655;
  initial
    n6656 = 1'b0;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6657 = clkena ? n5971 : current_privilege_level;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk or posedge n5967)
    if (n5967)
      n6658 <= 3'b000;
    else
      n6658 <= n6657;
  /* TG68K_FPU.vhd:3633:9  */
  assign n6661 = ~n5967;
  /* TG68K_FPU.vhd:3633:9  */
  assign n6662 = clkena & n6661;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6663 = n6662 ? n6250 : cir_handshake_state;
  /* TG68K_FPU.vhd:3663:17  */
  always @(posedge clk)
    n6664 <= n6663;
  initial
    n6664 = 3'b000;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6677 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6678 = clkena & n6677;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6679 = n6678 ? n5536 : operation_word_cir;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6680 <= n6679;
  initial
    n6680 = 16'b0000000000000000;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6681 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6682 = clkena & n6681;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6683 = n6682 ? n5538 : command_address_cir;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6684 <= n6683;
  initial
    n6684 = 32'b00000000000000000000000000000000;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6685 = clkena ? n5699 : fpu_state;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6686 <= 4'b0000;
    else
      n6686 <= n6685;
  /* TG68K_FPU.vhd:3619:17  */
  assign n6687 = clkena ? n5959 : fpu_busy_internal;
  /* TG68K_FPU.vhd:3619:17  */
  always @(posedge clk or posedge n5953)
    if (n5953)
      n6688 <= 1'b0;
    else
      n6688 <= n6687;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6691 = clkena ? n5548 : fsave_frame_format_latched;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6692 <= 8'b01100000;
    else
      n6692 <= n6691;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6693 = clkena ? n5551 : fpu_just_reset;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6694 <= 1'b0;
    else
      n6694 <= n6693;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6695 = clkena ? n5553 : movem_register_list;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6696 <= 8'b00000000;
    else
      n6696 <= n6695;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6697 = clkena ? n5555 : movem_direction;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6698 <= 1'b0;
    else
      n6698 <= n6697;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6699 = clkena ? n5559 : timeout_counter;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6700 <= 8'b00000000;
    else
      n6700 <= n6699;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6701 = clkena ? n5561 : fsave_counter;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6702 <= 6'b000000;
    else
      n6702 <= n6701;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6703 = clkena ? n5563 : frestore_frame_format;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6704 <= 8'b00000000;
    else
      n6704 <= n6703;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6709 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6710 = clkena & n6709;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6711 = n6710 ? n5569 : frestore_fp_temp;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6712 <= n6711;
  /* TG68K_FPU.vhd:1042:17  */
  assign n6713 = clkena ? n297 : fpu_operation;
  /* TG68K_FPU.vhd:1042:17  */
  always @(posedge clk or posedge n294)
    if (n294)
      n6714 <= 7'b0000000;
    else
      n6714 <= n6713;
  /* TG68K_FPU.vhd:1042:17  */
  assign n6715 = clkena ? n299 : source_reg;
  /* TG68K_FPU.vhd:1042:17  */
  always @(posedge clk or posedge n294)
    if (n294)
      n6716 <= 3'b000;
    else
      n6716 <= n6715;
  /* TG68K_FPU.vhd:1042:17  */
  assign n6717 = clkena ? n301 : dest_reg;
  /* TG68K_FPU.vhd:1042:17  */
  always @(posedge clk or posedge n294)
    if (n294)
      n6718 <= 3'b000;
    else
      n6718 <= n6717;
  /* TG68K_FPU.vhd:1042:17  */
  assign n6719 = clkena ? n303 : data_format;
  /* TG68K_FPU.vhd:1042:17  */
  always @(posedge clk or posedge n294)
    if (n294)
      n6720 <= 3'b000;
    else
      n6720 <= n6719;
  /* TG68K_FPU.vhd:1042:17  */
  assign n6721 = clkena ? n305 : ea_mode;
  /* TG68K_FPU.vhd:1042:17  */
  always @(posedge clk or posedge n294)
    if (n294)
      n6722 <= 3'b000;
    else
      n6722 <= n6721;
  /* TG68K_FPU.vhd:1042:17  */
  assign n6723 = clkena ? n307 : ea_register;
  /* TG68K_FPU.vhd:1042:17  */
  always @(posedge clk or posedge n294)
    if (n294)
      n6724 <= 3'b000;
    else
      n6724 <= n6723;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6728 = clkena ? n5681 : exception_code_internal;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6729 <= 8'b00000000;
    else
      n6729 <= n6728;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6730 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6731 = clkena & n6730;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6732 = n6731 ? n5574 : alu_start_operation;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6733 <= n6732;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6734 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6735 = clkena & n6734;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6736 = n6735 ? n5576 : alu_operation_code;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6737 <= n6736;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6738 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6739 = clkena & n6738;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6740 = n6739 ? n5578 : alu_operand_a;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6741 <= n6740;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6742 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6743 = clkena & n6742;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6744 = n6743 ? n5580 : alu_operand_b;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6745 <= n6744;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6746 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6747 = clkena & n6746;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6748 = n6747 ? n5583 : trans_start_operation;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6749 <= n6748;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6750 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6751 = clkena & n6750;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6752 = n6751 ? n5585 : trans_operation_code;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6753 <= n6752;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6754 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6755 = clkena & n6754;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6756 = n6755 ? n5587 : trans_operand;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6757 <= n6756;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6758 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6759 = clkena & n6758;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6760 = n6759 ? n5589 : final_result;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6761 <= n6760;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6762 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6763 = clkena & n6762;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6764 = n6763 ? n5591 : final_overflow;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6765 <= n6764;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6766 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6767 = clkena & n6766;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6768 = n6767 ? n5593 : final_underflow;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6769 <= n6768;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6770 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6771 = clkena & n6770;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6772 = n6771 ? n5595 : final_inexact;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6773 <= n6772;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6774 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6775 = clkena & n6774;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6776 = n6775 ? n5597 : final_invalid;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6777 <= n6776;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6778 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6779 = clkena & n6778;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6780 = n6779 ? n5599 : result_data;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6781 <= n6780;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6783 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6784 = clkena & n6783;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6785 = n6784 ? n5601 : converter_start;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6786 <= n6785;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6787 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6788 = clkena & n6787;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6789 = n6788 ? n5603 : converter_source_format;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6790 <= n6789;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6791 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6792 = clkena & n6791;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6793 = n6792 ? n5605 : converter_dest_format;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6794 <= n6793;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6795 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6796 = clkena & n6795;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6797 = n6796 ? n5607 : converter_data_in;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6798 <= n6797;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6799 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6800 = clkena & n6799;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6801 = n6800 ? n5609 : rom_offset;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6802 <= n6801;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6803 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6804 = clkena & n6803;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6805 = n6804 ? n5611 : rom_read_enable;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6806 <= n6805;
  /* TG68K_FPU.vhd:1179:9  */
  always @(n743)
    n6807 <= 1'b0;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6808 = clkena ? n5613 : movem_predecrement;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6809 <= 1'b0;
    else
      n6809 <= n6808;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6810 = clkena ? n5615 : movem_postincrement;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6811 <= 1'b0;
    else
      n6811 <= n6810;
  /* TG68K_FPU.vhd:3580:9  */
  assign n6812 = ~n5934;
  /* TG68K_FPU.vhd:3580:9  */
  assign n6813 = clkena & n6812;
  /* TG68K_FPU.vhd:3585:17  */
  assign n6814 = n6813 ? n5944 : movem_reg_data_in;
  /* TG68K_FPU.vhd:3585:17  */
  always @(posedge clk)
    n6815 <= n6814;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6832 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6833 = clkena & n6832;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6834 = n6833 ? n5623 : fp_to_int_shift;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6835 <= n6834;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6836 = ~n743;
  /* TG68K_FPU.vhd:1179:9  */
  assign n6837 = clkena & n6836;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6838 = n6837 ? n5625 : fp_to_int_result;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk)
    n6839 <= n6838;
  /* TG68K_FPU.vhd:1230:17  */
  assign n6840 = clkena ? n5337 : n6841;
  /* TG68K_FPU.vhd:1230:17  */
  always @(posedge clk or posedge n743)
    if (n743)
      n6841 <= 32'b00000000000000000000000000000000;
    else
      n6841 <= n6840;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6842 = n752[2]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6843 = ~n6842;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6844 = n752[1]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6845 = ~n6844;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6846 = n6843 & n6845;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6847 = n6843 & n6844;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6848 = n6842 & n6845;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6849 = n6842 & n6844;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6850 = n752[0]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6851 = ~n6850;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6852 = n6846 & n6851;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6853 = n6846 & n6850;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6854 = n6847 & n6851;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6855 = n6847 & n6850;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6856 = n6848 & n6851;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6857 = n6848 & n6850;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6858 = n6849 & n6851;
  /* TG68K_FPU.vhd:1236:49  */
  assign n6859 = n6849 & n6850;
  assign n6860 = fp_registers[79:0]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6861 = n6852 ? fp_reg_write_data : n6860;
  assign n6862 = fp_registers[159:80]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6863 = n6853 ? fp_reg_write_data : n6862;
  assign n6864 = fp_registers[239:160]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6865 = n6854 ? fp_reg_write_data : n6864;
  assign n6866 = fp_registers[319:240]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6867 = n6855 ? fp_reg_write_data : n6866;
  assign n6868 = fp_registers[399:320]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6869 = n6856 ? fp_reg_write_data : n6868;
  assign n6870 = fp_registers[479:400]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6871 = n6857 ? fp_reg_write_data : n6870;
  assign n6872 = fp_registers[559:480]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6873 = n6858 ? fp_reg_write_data : n6872;
  assign n6874 = fp_registers[639:560]; // extract
  /* TG68K_FPU.vhd:1236:49  */
  assign n6875 = n6859 ? fp_reg_write_data : n6874;
  assign n6876 = {n6875, n6873, n6871, n6869, n6867, n6865, n6863, n6861};
  /* TG68K_FPU.vhd:1510:113  */
  assign n6878 = {7'b0, n1279};  //  uext
  /* TG68K_FPU.vhd:1510:113  */
  assign n6879 = n6878 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1510:113  */
  assign n6880 = fp_registers[639:79]; // extract
  assign n6882 = {79'bX, n6880};
  /* TG68K_FPU.vhd:1525:111  */
  assign n6883 = n6882[n1310 * 80 +: 80]; //(Bmux)
  assign n6884 = n6883[0]; // extract
  /* TG68K_FPU.vhd:1526:126  */
  assign n6886 = {7'b0, n1316};  //  uext
  /* TG68K_FPU.vhd:1526:126  */
  assign n6887 = n6886 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1541:107  */
  assign n6888 = fp_registers[n1346 * 80 +: 80]; //(Bmux)
  /* TG68K_FPU.vhd:1578:101  */
  assign n6889 = fp_registers[n1438 * 80 +: 80]; //(Bmux)
  /* TG68K_FPU.vhd:1578:100  */
  assign n6890 = fp_registers[639:79]; // extract
  /* TG68K_FPU.vhd:1541:107  */
  assign n6892 = {79'bX, n6890};
  /* TG68K_FPU.vhd:1905:102  */
  assign n6893 = n6892[n1980 * 80 +: 80]; //(Bmux)
  assign n6894 = n6893[0]; // extract
  /* TG68K_FPU.vhd:1906:118  */
  assign n6896 = {7'b0, n1985};  //  uext
  /* TG68K_FPU.vhd:1906:118  */
  assign n6897 = n6896 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1907:118  */
  assign n6899 = {7'b0, n1993};  //  uext
  /* TG68K_FPU.vhd:1907:118  */
  assign n6900 = n6899 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1907:118  */
  assign n6901 = fp_registers[639:79]; // extract
  assign n6903 = {79'bX, n6901};
  /* TG68K_FPU.vhd:1916:102  */
  assign n6904 = n6903[n2001 * 80 +: 80]; //(Bmux)
  assign n6905 = n6904[0]; // extract
  /* TG68K_FPU.vhd:1916:143  */
  assign n6906 = fp_registers[639:65]; // extract
  assign n6908 = {65'bX, n6906};
  /* TG68K_FPU.vhd:1917:118  */
  assign n6909 = n6908[n2006 * 80 +: 80]; //(Bmux)
  assign n6910 = n6909[9:0]; // extract
  /* TG68K_FPU.vhd:1917:159  */
  assign n6911 = fp_registers[639:44]; // extract
  assign n6913 = {44'bX, n6911};
  /* TG68K_FPU.vhd:1918:118  */
  assign n6914 = n6913[n2014 * 80 +: 80]; //(Bmux)
  assign n6915 = n6914[19:0]; // extract
  /* TG68K_FPU.vhd:1933:89  */
  assign n6917 = {7'b0, n2037};  //  uext
  /* TG68K_FPU.vhd:1933:89  */
  assign n6918 = n6917 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1936:92  */
  assign n6920 = {7'b0, n2044};  //  uext
  /* TG68K_FPU.vhd:1936:92  */
  assign n6921 = n6920 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1936:92  */
  assign n6922 = fp_registers[639:79]; // extract
  assign n6924 = {79'bX, n6922};
  /* TG68K_FPU.vhd:1938:97  */
  assign n6925 = n6924[n2051 * 80 +: 80]; //(Bmux)
  assign n6926 = n6925[0]; // extract
  /* TG68K_FPU.vhd:1947:117  */
  assign n6928 = {7'b0, n2059};  //  uext
  /* TG68K_FPU.vhd:1947:117  */
  assign n6929 = n6928 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1950:120  */
  assign n6931 = {7'b0, n2068};  //  uext
  /* TG68K_FPU.vhd:1950:120  */
  assign n6932 = n6931 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1950:120  */
  assign n6933 = fp_registers[639:79]; // extract
  assign n6935 = {79'bX, n6933};
  /* TG68K_FPU.vhd:1952:105  */
  assign n6936 = n6935[n2077 * 80 +: 80]; //(Bmux)
  assign n6937 = n6936[0]; // extract
  /* TG68K_FPU.vhd:1960:125  */
  assign n6939 = {7'b0, n2085};  //  uext
  /* TG68K_FPU.vhd:1960:125  */
  assign n6940 = n6939 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1963:128  */
  assign n6942 = {7'b0, n2094};  //  uext
  /* TG68K_FPU.vhd:1963:128  */
  assign n6943 = n6942 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1968:155  */
  assign n6945 = {7'b0, n2103};  //  uext
  /* TG68K_FPU.vhd:1968:155  */
  assign n6946 = n6945 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1978:146  */
  assign n6948 = {7'b0, n2122};  //  uext
  /* TG68K_FPU.vhd:1978:146  */
  assign n6949 = n6948 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1981:184  */
  assign n6951 = {7'b0, n2129};  //  uext
  /* TG68K_FPU.vhd:1981:184  */
  assign n6952 = n6951 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:1981:184  */
  assign n6953 = fp_registers[639:79]; // extract
  /* TG68K_FPU.vhd:1230:17  */
  assign n6955 = {79'bX, n6953};
  /* TG68K_FPU.vhd:1991:105  */
  assign n6956 = n6955[n2147 * 80 +: 80]; //(Bmux)
  /* TG68K_FPU.vhd:1179:9  */
  assign n6957 = n6956[0]; // extract
  /* TG68K_FPU.vhd:2006:120  */
  assign n6958 = fp_registers[n2172 * 80 +: 80]; //(Bmux)
  /* TG68K_FPU.vhd:2014:120  */
  assign n6959 = fp_registers[n2180 * 80 +: 80]; //(Bmux)
  /* TG68K_FPU.vhd:2180:87  */
  assign n6960 = fp_registers[n2922 * 80 +: 80]; //(Bmux)
  /* TG68K_FPU.vhd:3075:127  */
  assign n6962 = {7'b0, n4489};  //  uext
  /* TG68K_FPU.vhd:3075:127  */
  assign n6963 = n6962 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:3082:127  */
  assign n6965 = {7'b0, n4506};  //  uext
  /* TG68K_FPU.vhd:3082:127  */
  assign n6966 = n6965 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:3090:141  */
  assign n6967 = fp_registers[n4523 * 80 +: 80]; //(Bmux)
  assign n6968 = n6967[15:0]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6969 = n4878[2]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6970 = ~n6969;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6971 = n4878[1]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6972 = ~n6971;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6973 = n6970 & n6972;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6974 = n6970 & n6971;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6975 = n6969 & n6972;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6976 = n6969 & n6971;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6977 = n4878[0]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6978 = ~n6977;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6979 = n6973 & n6978;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6980 = n6973 & n6977;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6981 = n6974 & n6978;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6982 = n6974 & n6977;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6983 = n6975 & n6978;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6984 = n6975 & n6977;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6985 = n6976 & n6978;
  /* TG68K_FPU.vhd:3295:105  */
  assign n6986 = n6976 & n6977;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6987 = frestore_fp_temp[47:0]; // extract
  /* TG68K_FPU.vhd:3663:17  */
  assign n6988 = frestore_fp_temp[79:48]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6989 = n6979 ? frestore_data_in : n6988;
  /* TG68K_FPU.vhd:3633:9  */
  assign n6990 = frestore_fp_temp[127:80]; // extract
  /* TG68K_FPU.vhd:3663:17  */
  assign n6991 = frestore_fp_temp[159:128]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6992 = n6980 ? frestore_data_in : n6991;
  /* TG68K_FPU.vhd:3633:9  */
  assign n6993 = frestore_fp_temp[207:160]; // extract
  /* TG68K_FPU.vhd:3633:9  */
  assign n6994 = frestore_fp_temp[239:208]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6995 = n6981 ? frestore_data_in : n6994;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6996 = frestore_fp_temp[287:240]; // extract
  /* TG68K_FPU.vhd:3663:17  */
  assign n6997 = frestore_fp_temp[319:288]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n6998 = n6982 ? frestore_data_in : n6997;
  /* TG68K_FPU.vhd:3663:17  */
  assign n6999 = frestore_fp_temp[367:320]; // extract
  /* TG68K_FPU.vhd:3663:17  */
  assign n7000 = frestore_fp_temp[399:368]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n7001 = n6983 ? frestore_data_in : n7000;
  /* TG68K_FPU.vhd:3663:17  */
  assign n7002 = frestore_fp_temp[447:400]; // extract
  /* TG68K_FPU.vhd:3663:17  */
  assign n7003 = frestore_fp_temp[479:448]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n7004 = n6984 ? frestore_data_in : n7003;
  /* TG68K_FPU.vhd:3663:17  */
  assign n7005 = frestore_fp_temp[527:480]; // extract
  /* TG68K_FPU.vhd:3663:17  */
  assign n7006 = frestore_fp_temp[559:528]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n7007 = n6985 ? frestore_data_in : n7006;
  /* TG68K_FPU.vhd:3663:17  */
  assign n7008 = frestore_fp_temp[607:560]; // extract
  /* TG68K_FPU.vhd:1230:17  */
  assign n7009 = frestore_fp_temp[639:608]; // extract
  /* TG68K_FPU.vhd:3295:105  */
  assign n7010 = n6986 ? frestore_data_in : n7009;
  /* TG68K_FPU.vhd:1179:9  */
  assign n7011 = {n7010, n7008, n7007, n7005, n7004, n7002, n7001, n6999, n6998, n6996, n6995, n6993, n6992, n6990, n6989, n6987};
  /* TG68K_FPU.vhd:3301:105  */
  assign n7012 = n4895[2]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7013 = ~n7012;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7014 = n4895[1]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7015 = ~n7014;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7016 = n7013 & n7015;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7017 = n7013 & n7014;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7018 = n7012 & n7015;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7019 = n7012 & n7014;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7020 = n4895[0]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7021 = ~n7020;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7022 = n7016 & n7021;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7023 = n7016 & n7020;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7024 = n7017 & n7021;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7025 = n7017 & n7020;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7026 = n7018 & n7021;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7027 = n7018 & n7020;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7028 = n7019 & n7021;
  /* TG68K_FPU.vhd:3301:105  */
  assign n7029 = n7019 & n7020;
  /* TG68K_FPU.vhd:1066:9  */
  assign n7030 = frestore_fp_temp[15:0]; // extract
  /* TG68K_FPU.vhd:1230:17  */
  assign n7031 = frestore_fp_temp[47:16]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7032 = n7022 ? frestore_data_in : n7031;
  /* TG68K_FPU.vhd:1230:17  */
  assign n7033 = frestore_fp_temp[95:48]; // extract
  /* TG68K_FPU.vhd:1230:17  */
  assign n7034 = frestore_fp_temp[127:96]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7035 = n7023 ? frestore_data_in : n7034;
  /* TG68K_FPU.vhd:1230:17  */
  assign n7036 = frestore_fp_temp[175:128]; // extract
  assign n7037 = frestore_fp_temp[207:176]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7038 = n7024 ? frestore_data_in : n7037;
  /* TG68K_FPU.vhd:4100:17  */
  assign n7039 = frestore_fp_temp[255:208]; // extract
  /* TG68K_FPU.vhd:4100:17  */
  assign n7040 = frestore_fp_temp[287:256]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7041 = n7025 ? frestore_data_in : n7040;
  /* TG68K_FPU.vhd:4100:17  */
  assign n7042 = frestore_fp_temp[335:288]; // extract
  assign n7043 = frestore_fp_temp[367:336]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7044 = n7026 ? frestore_data_in : n7043;
  assign n7045 = frestore_fp_temp[415:368]; // extract
  /* TG68K_FPU.vhd:4100:17  */
  assign n7046 = frestore_fp_temp[447:416]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7047 = n7027 ? frestore_data_in : n7046;
  /* TG68K_FPU.vhd:4103:33  */
  assign n7048 = frestore_fp_temp[495:448]; // extract
  assign n7049 = frestore_fp_temp[527:496]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7050 = n7028 ? frestore_data_in : n7049;
  /* TG68K_FPU.vhd:4103:33  */
  assign n7051 = frestore_fp_temp[575:528]; // extract
  assign n7052 = frestore_fp_temp[607:576]; // extract
  /* TG68K_FPU.vhd:3301:105  */
  assign n7053 = n7029 ? frestore_data_in : n7052;
  assign n7054 = frestore_fp_temp[639:608]; // extract
  /* TG68K_FPU.vhd:4131:41  */
  assign n7055 = {n7054, n7053, n7051, n7050, n7048, n7047, n7045, n7044, n7042, n7041, n7039, n7038, n7036, n7035, n7033, n7032, n7030};
  /* TG68K_FPU.vhd:3307:105  */
  assign n7056 = n4912[2]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7057 = ~n7056;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7058 = n4912[1]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7059 = ~n7058;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7060 = n7057 & n7059;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7061 = n7057 & n7058;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7062 = n7056 & n7059;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7063 = n7056 & n7058;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7064 = n4912[0]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7065 = ~n7064;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7066 = n7060 & n7065;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7067 = n7060 & n7064;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7068 = n7061 & n7065;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7069 = n7061 & n7064;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7070 = n7062 & n7065;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7071 = n7062 & n7064;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7072 = n7063 & n7065;
  /* TG68K_FPU.vhd:3307:105  */
  assign n7073 = n7063 & n7064;
  /* TG68K_FPU.vhd:4110:41  */
  assign n7074 = frestore_fp_temp[15:0]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7075 = n7066 ? n4914 : n7074;
  /* TG68K_FPU.vhd:4111:49  */
  assign n7076 = frestore_fp_temp[79:16]; // extract
  assign n7077 = frestore_fp_temp[95:80]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7078 = n7067 ? n4914 : n7077;
  assign n7079 = frestore_fp_temp[159:96]; // extract
  assign n7080 = frestore_fp_temp[175:160]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7081 = n7068 ? n4914 : n7080;
  assign n7082 = frestore_fp_temp[239:176]; // extract
  /* TG68K_FPU.vhd:4105:49  */
  assign n7083 = frestore_fp_temp[255:240]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7084 = n7069 ? n4914 : n7083;
  /* TG68K_FPU.vhd:4105:49  */
  assign n7085 = frestore_fp_temp[319:256]; // extract
  assign n7086 = frestore_fp_temp[335:320]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7087 = n7070 ? n4914 : n7086;
  /* TG68K_FPU.vhd:4105:84  */
  assign n7088 = frestore_fp_temp[399:336]; // extract
  assign n7089 = frestore_fp_temp[415:400]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7090 = n7071 ? n4914 : n7089;
  /* TG68K_FPU.vhd:4097:27  */
  assign n7091 = frestore_fp_temp[479:416]; // extract
  /* TG68K_FPU.vhd:4093:9  */
  assign n7092 = frestore_fp_temp[495:480]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7093 = n7072 ? n4914 : n7092;
  assign n7094 = frestore_fp_temp[559:496]; // extract
  /* TG68K_FPU.vhd:4094:26  */
  assign n7095 = frestore_fp_temp[575:560]; // extract
  /* TG68K_FPU.vhd:3307:105  */
  assign n7096 = n7073 ? n4914 : n7095;
  assign n7097 = frestore_fp_temp[639:576]; // extract
  assign n7098 = {n7097, n7096, n7094, n7093, n7091, n7090, n7088, n7087, n7085, n7084, n7082, n7081, n7079, n7078, n7076, n7075};
  /* TG68K_FPU.vhd:3310:157  */
  assign n7100 = {7'b0, n4926};  //  uext
  /* TG68K_FPU.vhd:3310:157  */
  assign n7101 = n7100 * 10'b0001010000; // umul
  /* TG68K_FPU.vhd:3589:75  */
  assign n7102 = fp_registers[n5940 * 80 +: 80]; //(Bmux)
endmodule

