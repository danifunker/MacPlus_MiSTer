///////////////////////////////////////////////////////////////////////////////
// Title      : VIA 6522
///////////////////////////////////////////////////////////////////////////////
// Author     : Gideon Zweijtzer  <gideon.zweijtzer@gmail.com>
///////////////////////////////////////////////////////////////////////////////
// Description: This module implements the 6522 VIA chip.
//              A LOT OF REVERSE ENGINEERING has been done to make this module
//              as accurate as it is now. Thanks to gyurco for ironing out some
//              differences that were left unnoticed.
///////////////////////////////////////////////////////////////////////////////
// License:     GPL 3.0 - Free to use, distribute and change to your own needs.
//              Leaving a reference to the author will be highly appreciated.
///////////////////////////////////////////////////////////////////////////////

module via6522 (
    input  wire        clock,
    input  wire        rising,
    input  wire        falling,
    input  wire        reset,
    
    input  wire [3:0]  addr,
    input  wire        wen,
    input  wire        ren,
    input  wire [7:0]  data_in,
    output reg  [7:0]  data_out,

    output reg         phi2_ref,

    // pio
    output wire [7:0]  port_a_o,
    output wire [7:0]  port_a_t,
    input  wire [7:0]  port_a_i,
    
    output wire [7:0]  port_b_o,
    output wire [7:0]  port_b_t,
    input  wire [7:0]  port_b_i,

    // handshake pins
    input  wire        ca1_i,

    output wire        ca2_o,
    input  wire        ca2_i,
    output wire        ca2_t,
    
    output wire        cb1_o,
    input  wire        cb1_i,
    output wire        cb1_t,
    
    output wire        cb2_o,
    input  wire        cb2_i,
    output wire        cb2_t,

    output wire        irq
);

    localparam [15:0] latch_reset_pattern = 16'h5550;

    // PIO signals (replaces record type)
    reg [7:0] pio_i_pra  = 8'h00;
    reg [7:0] pio_i_ddra = 8'h00;
    reg [7:0] pio_i_prb  = 8'h00;
    reg [7:0] pio_i_ddrb = 8'h00;
    
    reg [7:0] port_a_c = 8'h00;
    reg [7:0] port_b_c = 8'h00;
    
    reg [6:0] irq_mask   = 7'h00;
    reg [6:0] irq_flags  = 7'h00;
    reg [6:0] irq_events = 7'h00;
    reg       irq_out;
    
    reg [15:0] timer_a_latch = latch_reset_pattern;
    reg [15:0] timer_b_latch = latch_reset_pattern;
    reg [15:0] timer_a_count = latch_reset_pattern;
    reg [15:0] timer_b_count = latch_reset_pattern;
    reg        timer_a_out;
    reg        timer_b_tick;
                         
    reg [7:0] acr = 8'h00;
    reg [7:0] pcr = 8'h00;
    reg [7:0] shift_reg = 8'h00;
    reg       serport_en;
    reg       ser_cb2_o;
    reg       hs_cb2_o;
    reg       cb1_t_int;
    reg       cb1_o_int;
    reg       cb2_t_int;
    reg       cb2_o_int;

    // Aliases for irq_events
    wire ca2_event     = irq_events[0];
    wire ca1_event     = irq_events[1];
    wire serial_event  = irq_events[2];
    wire cb2_event     = irq_events[3];
    wire cb1_event     = irq_events[4];
    wire timer_b_event = irq_events[5];
    wire timer_a_event = irq_events[6];

    // Aliases for irq_flags
    wire ca2_flag     = irq_flags[0];
    wire ca1_flag     = irq_flags[1];
    wire serial_flag  = irq_flags[2];
    wire cb2_flag     = irq_flags[3];
    wire cb1_flag     = irq_flags[4];
    wire timer_b_flag = irq_flags[5];
    wire timer_a_flag = irq_flags[6];

    // Aliases for ACR bits
    wire       tmr_a_output_en       = acr[7];
    wire       tmr_a_freerun         = acr[6];
    wire       tmr_b_count_mode      = acr[5];
    wire       shift_dir             = acr[4];
    wire [1:0] shift_clk_sel         = acr[3:2];
    wire [2:0] shift_mode_control    = acr[4:2];
    wire       pb_latch_en           = acr[1];
    wire       pa_latch_en           = acr[0];
    
    // Aliases for PCR bits
    wire       cb2_is_output         = pcr[7];
    wire       cb2_edge_select       = pcr[6];
    wire       cb2_no_irq_clr        = pcr[5];
    wire [1:0] cb2_out_mode          = pcr[6:5];
    wire       cb1_edge_select       = pcr[4];
    
    wire       ca2_is_output         = pcr[3];
    wire       ca2_edge_select       = pcr[2];
    wire       ca2_no_irq_clr        = pcr[1];
    wire [1:0] ca2_out_mode          = pcr[2:1];
    wire       ca1_edge_select       = pcr[0];
    
    reg [7:0] ira = 8'h00;
    reg [7:0] irb = 8'h00;

    reg write_t1c_l;
    reg write_t1c_h;
    reg write_t2c_h;

    reg ca1_c = 1'b0;
    reg ca2_c = 1'b0;
    reg cb1_c = 1'b0;
    reg cb2_c = 1'b0;
    reg ca1_d = 1'b0;
    reg ca2_d = 1'b0;
    reg cb1_d = 1'b0;
    reg cb2_d = 1'b0;
    
    reg ca2_handshake_o = 1'b1;
    reg ca2_pulse_o = 1'b1;
    reg cb2_handshake_o = 1'b1;
    reg cb2_pulse_o = 1'b1;
    reg shift_active;

    // Assignments
    assign irq = irq_out;
    
    always @(*) begin
        write_t1c_l = ((addr == 4'h4 || addr == 4'h6) && wen && falling);
        write_t1c_h = (addr == 4'h5 && wen && falling);
        write_t2c_h = (addr == 4'h9 && wen && falling);
    end

    always @(*) begin
        irq_events[1] = (ca1_c ^ ca1_d) & (ca1_d ^ ca1_edge_select);
        irq_events[0] = (ca2_c ^ ca2_d) & (ca2_d ^ ca2_edge_select);
        irq_events[4] = (cb1_c ^ cb1_d) & (cb1_d ^ cb1_edge_select);
        irq_events[3] = (cb2_c ^ cb2_d) & (cb2_d ^ cb2_edge_select);
    end

    assign ca2_t = ca2_is_output;
    
    always @(*) begin
        cb2_t_int = serport_en ? shift_dir : cb2_is_output;
        cb2_o_int = serport_en ? ser_cb2_o : hs_cb2_o;
    end

    assign cb1_t = cb1_t_int;
    assign cb1_o = cb1_o_int;
    assign cb2_t = cb2_t_int;
    assign cb2_o = cb2_o_int;

    assign ca2_o = (ca2_out_mode == 2'b00) ? ca2_handshake_o :
                   (ca2_out_mode == 2'b01) ? ca2_pulse_o :
                   (ca2_out_mode == 2'b10) ? 1'b0 : 1'b1;
        
    always @(*) begin
        hs_cb2_o = (cb2_out_mode == 2'b00) ? cb2_handshake_o :
                   (cb2_out_mode == 2'b01) ? cb2_pulse_o :
                   (cb2_out_mode == 2'b10) ? 1'b0 : 1'b1;
    end

    always @(*) begin
        if ((irq_flags & irq_mask) == 7'h00) begin
            irq_out = 1'b0;
        end else begin
            irq_out = 1'b1;
        end
    end

    always @(posedge clock) begin
        if (rising) begin
            phi2_ref <= 1'b1;
        end else if (falling) begin
            phi2_ref <= 1'b0;
        end
    end

    always @(posedge clock) begin
        // CA1/CA2/CB1/CB2 edge detect flipflops
        ca1_c <= ca1_i;
        ca2_c <= ca2_i;
        if (cb1_t_int == 1'b0) begin
            cb1_c <= cb1_i;
        end else begin
            cb1_c <= cb1_o_int;
        end
        if (cb2_t_int == 1'b0) begin
            cb2_c <= cb2_i;
        end else begin
            cb2_c <= cb2_o_int;
        end

        ca1_d <= ca1_c;
        ca2_d <= ca2_c;
        cb1_d <= cb1_c;
        cb2_d <= cb2_c;

        // input registers
        port_a_c <= port_a_i;
        port_b_c <= port_b_i;

        // input latch emulation
        if (pa_latch_en == 1'b0 || ca1_event == 1'b1) begin
            ira <= port_a_c;
        end
        
        if (pb_latch_en == 1'b0 || cb1_event == 1'b1) begin
            irb <= port_b_c;
        end

        // CA2 logic
        if (ca1_event == 1'b1) begin
            ca2_handshake_o <= 1'b1;
        end else if ((ren == 1'b1 || wen == 1'b1) && addr == 4'h1 && falling == 1'b1) begin
            ca2_handshake_o <= 1'b0;
        end
        
        if (falling == 1'b1) begin
            if ((ren == 1'b1 || wen == 1'b1) && addr == 4'h1) begin
                ca2_pulse_o <= 1'b0;
            end else begin
                ca2_pulse_o <= 1'b1;
            end
        end

        // CB2 logic
        if (cb1_event == 1'b1) begin
            cb2_handshake_o <= 1'b1;
        end else if ((ren == 1'b1 || wen == 1'b1) && addr == 4'h0 && falling == 1'b1) begin
            cb2_handshake_o <= 1'b0;
        end
        
        if (falling == 1'b1) begin
            if ((ren == 1'b1 || wen == 1'b1) && addr == 4'h0) begin
                cb2_pulse_o <= 1'b0;
            end else begin
                cb2_pulse_o <= 1'b1;
            end
        end

        // Interrupt logic
        irq_flags <= irq_flags | irq_events;

        // Writes
        if (wen == 1'b1 && falling == 1'b1) begin
            case (addr)
                4'h0: begin // ORB
                    pio_i_prb <= data_in;
                    if (cb2_no_irq_clr == 1'b0) begin
                        irq_flags[3] <= 1'b0;
                    end
                    irq_flags[4] <= 1'b0;
                end
                
                4'h1: begin // ORA
                    pio_i_pra <= data_in;
                    if (ca2_no_irq_clr == 1'b0) begin
                        irq_flags[0] <= 1'b0;
                    end
                    irq_flags[1] <= 1'b0;
                end
                    
                4'h2: begin // DDRB
                    pio_i_ddrb <= data_in;
                end
                
                4'h3: begin // DDRA
                    pio_i_ddra <= data_in;
                end
                    
                4'h4: begin // TA LO counter (write=latch)
                    timer_a_latch[7:0] <= data_in;
                end
                    
                4'h5: begin // TA HI counter
                    timer_a_latch[15:8] <= data_in;
                    irq_flags[6] <= 1'b0;
                end
                    
                4'h6: begin // TA LO latch
                    timer_a_latch[7:0] <= data_in;
                end
                    
                4'h7: begin // TA HI latch
                    timer_a_latch[15:8] <= data_in;
                    irq_flags[6] <= 1'b0;
                end
                    
                4'h8: begin // TB LO latch
                    timer_b_latch[7:0] <= data_in;
                end
                    
                4'h9: begin // TB HI counter
                    irq_flags[5] <= 1'b0;
                end
                    
                4'hA: begin // Serial port
                    irq_flags[2] <= 1'b0;
                end
                    
                4'hB: begin // ACR (Auxiliary Control Register)
                    acr <= data_in;
                end
                    
                4'hC: begin // PCR (Peripheral Control Register)
                    pcr <= data_in;
                end
                                    
                4'hD: begin // IFR
                    irq_flags <= irq_flags & ~data_in[6:0];
                end
                    
                4'hE: begin // IER
                    if (data_in[7] == 1'b1) begin // set
                        irq_mask <= irq_mask | data_in[6:0];
                    end else begin // clear
                        irq_mask <= irq_mask & ~data_in[6:0];
                    end
                end
                
                4'hF: begin // ORA no handshake
                    pio_i_pra <= data_in;
                end
                
                default: begin
                end
            endcase
        end
        
        // Reads - Output only
        data_out <= 8'h00;
        case (addr)
            4'h0: begin // ORB
                // Port B reads its own output register for pins set to output.
                data_out <= (pio_i_prb & pio_i_ddrb) | (irb & ~pio_i_ddrb);
                if (tmr_a_output_en == 1'b1) begin
                    data_out[7] <= timer_a_out;
                end
            end
            4'h1: begin // ORA
                data_out <= ira;
            end
            4'h2: begin // DDRB
                data_out <= pio_i_ddrb;
            end
            4'h3: begin // DDRA
                data_out <= pio_i_ddra;
            end
            4'h4: begin // TA LO counter
                data_out <= timer_a_count[7:0];
            end
            4'h5: begin // TA HI counter
                data_out <= timer_a_count[15:8];
            end
            4'h6: begin // TA LO latch
                data_out <= timer_a_latch[7:0];
            end
            4'h7: begin // TA HI latch
                data_out <= timer_a_latch[15:8];
            end
            4'h8: begin // TA LO counter
                data_out <= timer_b_count[7:0];
            end
            4'h9: begin // TA HI counter
                data_out <= timer_b_count[15:8];
            end
            4'hA: begin // SR
                data_out <= shift_reg;
            end
            4'hB: begin // ACR
                data_out <= acr;
            end
            4'hC: begin // PCR
                data_out <= pcr;
            end
            4'hD: begin // IFR
                data_out <= {irq_out, irq_flags};
            end
            4'hE: begin // IER
                data_out <= {1'b1, irq_mask};
            end
            4'hF: begin // ORA
                data_out <= ira;
            end
            default: begin
            end
        endcase
        
        // Read actions
        if (ren == 1'b1 && falling == 1'b1) begin
            case (addr)
                4'h0: begin // ORB
                    if (cb2_no_irq_clr == 1'b0) begin
                        irq_flags[3] <= 1'b0;
                    end
                    irq_flags[4] <= 1'b0;
                end
                                            
                4'h1: begin // ORA
                    if (ca2_no_irq_clr == 1'b0) begin
                        irq_flags[0] <= 1'b0;
                    end
                    irq_flags[1] <= 1'b0;
                end
                    
                4'h4: begin // TA LO counter
                    irq_flags[6] <= 1'b0;
                end
                    
                4'h8: begin // TB LO counter
                    irq_flags[5] <= 1'b0;
                end
                    
                4'hA: begin // SR
                    irq_flags[2] <= 1'b0;
                end
    
                default: begin
                end
            endcase
        end

        if (reset == 1'b1) begin
            pio_i_pra       <= 8'h00;
            pio_i_ddra      <= 8'h00;
            pio_i_prb       <= 8'h00;
            pio_i_ddrb      <= 8'h00;
            irq_mask        <= 7'h00;
            irq_flags       <= 7'h00;
            acr             <= 8'h00;
            pcr             <= 8'h00;
            ca2_handshake_o <= 1'b1;
            ca2_pulse_o     <= 1'b1;
            cb2_handshake_o <= 1'b1;
            cb2_pulse_o     <= 1'b1;
            timer_a_latch   <= latch_reset_pattern;
            timer_b_latch   <= latch_reset_pattern;
        end
    end

    // PIO Out select
    assign port_a_o = pio_i_pra;
    assign port_b_o[6:0] = pio_i_prb[6:0];
    assign port_b_o[7] = (tmr_a_output_en == 1'b0) ? pio_i_prb[7] : timer_a_out;
    
    assign port_a_t = pio_i_ddra;
    assign port_b_t[6:0] = pio_i_ddrb[6:0];
    assign port_b_t[7] = pio_i_ddrb[7] | tmr_a_output_en;

    // Timer A
    reg        timer_a_reload = 1'b0;
    reg        timer_a_toggle = 1'b1;
    reg        timer_a_may_interrupt = 1'b0;

    always @(posedge clock) begin
        if (falling == 1'b1) begin
            // always count, or load
                
            if (timer_a_reload == 1'b1) begin
                timer_a_count <= timer_a_latch;
                if (write_t1c_l == 1'b1) begin
                    timer_a_count[7:0] <= data_in;
                end
                timer_a_reload <= 1'b0;
                timer_a_may_interrupt <= timer_a_may_interrupt & tmr_a_freerun;
            end else begin
                if (timer_a_count == 16'h0000) begin
                    // generate an event if we were triggered
                    timer_a_reload <= 1'b1;
                end
                // Timer continues to count in both free run and one shot.
                timer_a_count <= timer_a_count - 16'h0001;
            end
        end
        
        if (rising == 1'b1) begin
            if (timer_a_event == 1'b1 && tmr_a_output_en == 1'b1) begin
                timer_a_toggle <= ~timer_a_toggle;
            end
        end

        if (write_t1c_h == 1'b1) begin
            timer_a_may_interrupt <= 1'b1;
            timer_a_toggle <= ~tmr_a_output_en;
            timer_a_count <= {data_in, timer_a_latch[7:0]};
            timer_a_reload <= 1'b0;
        end

        if (reset == 1'b1) begin
            timer_a_may_interrupt <= 1'b0;
            timer_a_toggle <= 1'b1;
            timer_a_count <= latch_reset_pattern;
            timer_a_reload <= 1'b0;
        end
    end

    assign timer_a_out = timer_a_toggle;
    assign timer_a_event = rising & timer_a_reload & timer_a_may_interrupt;

    // Timer B
    reg        timer_b_reload_lo = 1'b0;
    reg        timer_b_oneshot_trig = 1'b0;
    reg        timer_b_timeout = 1'b0;
    reg        pb6_c = 1'b0;
    reg        pb6_d = 1'b0;

    always @(posedge clock) begin
        reg timer_b_decrement;
        
        timer_b_decrement = 1'b0;

        if (rising == 1'b1) begin
            pb6_c <= port_b_i[6];
            pb6_d <= pb6_c;
        end
                        
        if (falling == 1'b1) begin
            timer_b_timeout <= 1'b0;
            timer_b_tick <= 1'b0;

            if (tmr_b_count_mode == 1'b1) begin
                if (pb6_d == 1'b1 && pb6_c == 1'b0) begin
                    timer_b_decrement = 1'b1;
                end
            end else begin // one shot or used for shift register
                timer_b_decrement = 1'b1;
            end
                
            if (timer_b_decrement == 1'b1) begin
                if (timer_b_count == 16'h0000) begin
                    if (timer_b_oneshot_trig == 1'b1) begin
                        timer_b_oneshot_trig <= 1'b0;
                        timer_b_timeout <= 1'b1;
                    end
                end
                if (timer_b_count[7:0] == 8'h00) begin
                    case (shift_mode_control)
                        3'b001, 3'b101, 3'b100: begin
                            timer_b_reload_lo <= 1'b1;
                            timer_b_tick <= 1'b1;
                        end
                        default: begin
                        end
                    endcase
                end
                timer_b_count <= timer_b_count - 16'h0001;
            end
            if (timer_b_reload_lo == 1'b1) begin
                timer_b_count[7:0] <= timer_b_latch[7:0];
                timer_b_reload_lo <= 1'b0;
            end
        end

        if (write_t2c_h == 1'b1) begin
            timer_b_count <= {data_in, timer_b_latch[7:0]};
            timer_b_oneshot_trig <= 1'b1;
        end

        if (reset == 1'b1) begin
            timer_b_count <= latch_reset_pattern;
            timer_b_reload_lo <= 1'b0;
            timer_b_oneshot_trig <= 1'b0;
        end
    end

    assign timer_b_event = rising & timer_b_timeout;

    // Serial port
    reg        trigger_serial;
    reg        shift_clock_d = 1'b1;
    reg        shift_clock = 1'b1;
    reg        shift_tick_r;
    reg        shift_tick_f;
    reg        shift_timer_tick;
    reg        ser_cb2_c = 1'b0;
    reg [2:0]  bit_cnt = 3'd0;
    reg        shift_pulse;

    always @(*) begin
        case (shift_clk_sel)
            2'b10: begin
                shift_pulse = 1'b1;
            end
                
            2'b00, 2'b01: begin
                shift_pulse = shift_timer_tick;
            end
            
            default: begin
                shift_pulse = shift_clock & ~shift_clock_d;
            end
        endcase

        if (shift_active == 1'b0) begin
            // Mode 0 still loads the shift register to external pulse (MMBEEB SD-Card interface uses this)
            if (shift_mode_control == 3'b000) begin
                shift_pulse = shift_clock & ~shift_clock_d;
            end else begin
                shift_pulse = 1'b0;
            end
        end
    end

    always @(posedge clock) begin
        ser_cb2_c <= cb2_i;

        if (rising == 1'b1) begin
            if (shift_active == 1'b0) begin
                if (shift_mode_control == 3'b000) begin
                    shift_clock <= cb1_i;
                end else begin
                    shift_clock <= 1'b1;
                end
            end else if (shift_clk_sel == 2'b11) begin
                shift_clock <= cb1_i;
            end else if (shift_pulse == 1'b1) begin
                shift_clock <= ~shift_clock;
            end

            shift_clock_d <= shift_clock;
        end

        if (falling == 1'b1) begin
            shift_timer_tick <= timer_b_tick;
        end

        if (reset == 1'b1) begin
            shift_clock <= 1'b1;
            shift_clock_d <= 1'b1;
        end
    end

    always @(*) begin
        cb1_t_int = (shift_clk_sel == 2'b11) ? 1'b0 : serport_en;
        cb1_o_int = shift_clock_d;
        ser_cb2_o = shift_reg[7];
    end

    always @(*) begin
        serport_en = shift_dir | shift_clk_sel[1] | shift_clk_sel[0];
        trigger_serial = ((ren == 1'b1 || wen == 1'b1) && addr == 4'hA);
        shift_tick_r = ~shift_clock_d & shift_clock;
        shift_tick_f = shift_clock_d & ~shift_clock;
    end

    always @(posedge clock) begin
        if (reset == 1'b1) begin
            shift_reg <= 8'hFF;
        end else if (falling == 1'b1) begin
            if (wen == 1'b1 && addr == 4'hA) begin
                shift_reg <= data_in;
            end else if (shift_dir == 1'b1 && shift_tick_f == 1'b1) begin // output
                shift_reg <= {shift_reg[6:0], shift_reg[7]};
            end else if (shift_dir == 1'b0 && shift_tick_r == 1'b1) begin // input
                shift_reg <= {shift_reg[6:0], ser_cb2_c};
            end
        end
    end

    // tell people that we're ready!
    assign serial_event = shift_tick_r & ~shift_active & rising & serport_en;

    always @(posedge clock) begin
        if (falling == 1'b1) begin
            if (shift_active == 1'b0 && shift_mode_control != 3'b000) begin
                if (trigger_serial == 1'b1) begin
                    bit_cnt <= 3'd7;
                    shift_active <= 1'b1;
                end
            end else begin // we're active
                if (shift_clk_sel == 2'b00) begin
                    shift_active <= shift_dir; // when '1' we're active, but for mode 000 we go inactive.
                end else if (shift_pulse == 1'b1 && shift_clock == 1'b1) begin
                    if (bit_cnt == 3'd0) begin
                        shift_active <= 1'b0;
                    end else begin
                        bit_cnt <= bit_cnt - 3'd1;
                    end
                end
            end
        end

        if (reset == 1'b1) begin
            shift_active <= 1'b0;
            bit_cnt <= 3'd0;
        end
    end

endmodule
