module TG68K_FPU_ConstantROM
  (input  clk,
   input  nReset,
   input  [6:0] rom_offset,
   input  read_enable,
   output [79:0] constant_out,
   output constant_valid);
  wire n3;
  wire n6;
  wire n8;
  wire n10;
  wire n12;
  wire n14;
  wire n16;
  wire n18;
  wire n20;
  wire n22;
  wire n24;
  wire n26;
  wire n28;
  wire n30;
  wire n32;
  wire n34;
  wire n36;
  wire n38;
  wire n40;
  wire n42;
  wire n44;
  wire n46;
  wire n48;
  wire [21:0] n49;
  reg [79:0] n73;
  wire n77;
  wire [79:0] n86;
  reg [79:0] n87;
  reg n88;
  assign constant_out = n87; //(module output)
  assign constant_valid = n88; //(module output)
  /* TG68K_FPU_ConstantROM.vhd:104:27  */
  assign n3 = ~nReset;
  /* TG68K_FPU_ConstantROM.vhd:112:41  */
  assign n6 = rom_offset == 7'b0000000;
  /* TG68K_FPU_ConstantROM.vhd:115:41  */
  assign n8 = rom_offset == 7'b0001011;
  /* TG68K_FPU_ConstantROM.vhd:118:41  */
  assign n10 = rom_offset == 7'b0001100;
  /* TG68K_FPU_ConstantROM.vhd:121:41  */
  assign n12 = rom_offset == 7'b0001101;
  /* TG68K_FPU_ConstantROM.vhd:124:41  */
  assign n14 = rom_offset == 7'b0001110;
  /* TG68K_FPU_ConstantROM.vhd:127:41  */
  assign n16 = rom_offset == 7'b0001111;
  /* TG68K_FPU_ConstantROM.vhd:130:41  */
  assign n18 = rom_offset == 7'b0110000;
  /* TG68K_FPU_ConstantROM.vhd:133:41  */
  assign n20 = rom_offset == 7'b0110001;
  /* TG68K_FPU_ConstantROM.vhd:136:41  */
  assign n22 = rom_offset == 7'b0110010;
  /* TG68K_FPU_ConstantROM.vhd:139:41  */
  assign n24 = rom_offset == 7'b0110011;
  /* TG68K_FPU_ConstantROM.vhd:142:41  */
  assign n26 = rom_offset == 7'b0110100;
  /* TG68K_FPU_ConstantROM.vhd:145:41  */
  assign n28 = rom_offset == 7'b0110101;
  /* TG68K_FPU_ConstantROM.vhd:148:41  */
  assign n30 = rom_offset == 7'b0110110;
  /* TG68K_FPU_ConstantROM.vhd:151:41  */
  assign n32 = rom_offset == 7'b0110111;
  /* TG68K_FPU_ConstantROM.vhd:154:41  */
  assign n34 = rom_offset == 7'b0111000;
  /* TG68K_FPU_ConstantROM.vhd:157:41  */
  assign n36 = rom_offset == 7'b0111001;
  /* TG68K_FPU_ConstantROM.vhd:160:41  */
  assign n38 = rom_offset == 7'b0111010;
  /* TG68K_FPU_ConstantROM.vhd:163:41  */
  assign n40 = rom_offset == 7'b0111011;
  /* TG68K_FPU_ConstantROM.vhd:166:41  */
  assign n42 = rom_offset == 7'b0111100;
  /* TG68K_FPU_ConstantROM.vhd:169:41  */
  assign n44 = rom_offset == 7'b0111101;
  /* TG68K_FPU_ConstantROM.vhd:172:41  */
  assign n46 = rom_offset == 7'b0111110;
  /* TG68K_FPU_ConstantROM.vhd:175:41  */
  assign n48 = rom_offset == 7'b0111111;
  assign n49 = {n48, n46, n44, n42, n40, n38, n36, n34, n32, n30, n28, n26, n24, n22, n20, n18, n16, n14, n12, n10, n8, n6};
  /* TG68K_FPU_ConstantROM.vhd:111:33  */
  always @*
    case (n49)
      22'b1000000000000000000000: n73 = 80'b01110101001001011100010001100000000100100111101010111100110010001111011010101111;
      22'b0100000000000000000000: n73 = 80'b01011010100100101001000101111111010101000111110101110011110010000000011100000001;
      22'b0010000000000000000000: n73 = 80'b01001101010010001100100101110110011101011000011010000001011101010000110000010111;
      22'b0001000000000000000000: n73 = 80'b01000110101000111100011000110011010000010101110101001100000111010010001110001101;
      22'b0000100000000000000000: n73 = 80'b01000011010100011010101001111110111010111111101110011101111110011101111010001110;
      22'b0000010000000000000000: n73 = 80'b01000001101010001001001110111010010001111100100110000000111010011000110011100000;
      22'b0000001000000000000000: n73 = 80'b01000000110100111000010011110000001111101001001111111111100111110100110110101010;
      22'b0000000100000000000000: n73 = 80'b01000000011010010011101110001011010110110101000001010110111000010110101100111100;
      22'b0000000010000000000000: n73 = 80'b01000000001101001000111000011011110010011011111100000100000000000000000000000000;
      22'b0000000001000000000000: n73 = 80'b01000000000110011011111010111100001000000000000000000000000000000000000000000000;
      22'b0000000000100000000000: n73 = 80'b01000000000011001001110001000000000000000000000000000000000000000000000000000000;
      22'b0000000000010000000000: n73 = 80'b01000000000001011100100000000000000000000000000000000000000000000000000000000000;
      22'b0000000000001000000000: n73 = 80'b01000000000000101010000000000000000000000000000000000000000000000000000000000000;
      22'b0000000000000100000000: n73 = 80'b00111111111111111000000000000000000000000000000000000000000000000000000000000000;
      22'b0000000000000010000000: n73 = 80'b01000000000000001001001101011101100011011101110110101010101010001010110000010111;
      22'b0000000000000001000000: n73 = 80'b00111111111111101011000101110010000101111111011111010001110011110111100110101100;
      22'b0000000000000000100000: n73 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
      22'b0000000000000000010000: n73 = 80'b00111111111111011101111001011011110110001010100100110111001010000111000110010101;
      22'b0000000000000000001000: n73 = 80'b00111111111111111011100010101010001110110010100101011100000101111111000010111100;
      22'b0000000000000000000100: n73 = 80'b01000000000000001010110111111000010101000101100010100010101110110100101010011010;
      22'b0000000000000000000010: n73 = 80'b00111111111111011001101000100000100110101000010011111011110011111111011110011000;
      22'b0000000000000000000001: n73 = 80'b01000000000000001100100100001111110110101010001000100001011010001100001000110101;
      default: n73 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* TG68K_FPU_ConstantROM.vhd:110:25  */
  assign n77 = read_enable ? 1'b1 : 1'b0;
  /* TG68K_FPU_ConstantROM.vhd:107:17  */
  assign n86 = read_enable ? n73 : n87;
  /* TG68K_FPU_ConstantROM.vhd:107:17  */
  always @(posedge clk or posedge n3)
    if (n3)
      n87 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n87 <= n86;
  /* TG68K_FPU_ConstantROM.vhd:107:17  */
  always @(posedge clk or posedge n3)
    if (n3)
      n88 <= 1'b0;
    else
      n88 <= n77;
endmodule

